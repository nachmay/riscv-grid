**** Created by MC2: Version 2013.12.00.f on 2025/06/23, 08:34:15 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  N16FF_SPSB_LEAFCELL
* Top Cell Name: LEAFCELL
* View Name:     schematic
* Netlisted on:  Jun  4 15:47:25 2014
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM


*.PIN vss
.SUBCKT ndio_mac PLUS MINUS 
.ends

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    BCELL_SD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_BCELL_SD TSMC_1 TSMC_2 VDDAI VDDI VSSI TSMC_3 
MM5 TSMC_2 TSMC_3 TSMC_4 VSSI nchpg_hcsr_mac l=20n nfin=2 m=1 
MM0 TSMC_1 TSMC_3 TSMC_5 VSSI nchpg_hcsr_mac l=20n nfin=2 m=1 
MM2 TSMC_4 TSMC_5 VSSI VSSI nchpd_hcsr_mac l=20n nfin=2 m=1 
MM1 TSMC_5 TSMC_4 VSSI VSSI nchpd_hcsr_mac l=20n nfin=2 m=1 
MM6 TSMC_5 TSMC_4 VDDAI VDDI pchpu_hcsr_mac l=20n nfin=1 m=1 
MM4 TSMC_4 TSMC_5 VDDAI VDDI pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_lvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_nand3_lvt_mac_pcell_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_lvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_lvt_mac_pcell_5
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_nor2_lvt_mac_pcell_5 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_6
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    XDRV_LA512_884_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_XDRV_LA512_884_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 VDDI VSSI TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 
MM37 TSMC_26 TSMC_30 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM36 TSMC_30 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM35 TSMC_22 TSMC_30 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM34 TSMC_30 TSMC_31 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM33 TSMC_31 TSMC_3 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MM21 TSMC_27 TSMC_33 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM16 TSMC_33 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM13 TSMC_23 TSMC_33 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM11 TSMC_33 TSMC_34 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM10 TSMC_34 TSMC_4 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MM3 TSMC_25 TSMC_35 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM2 TSMC_24 TSMC_36 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM23 TSMC_21 TSMC_35 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM20 TSMC_20 TSMC_36 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM28 TSMC_35 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM27 TSMC_36 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM26 TSMC_35 TSMC_37 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM18 TSMC_36 TSMC_38 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM12 TSMC_37 TSMC_2 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MP6 TSMC_38 TSMC_1 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MM39 TSMC_32 TSMC_9 VDDI VDDI pch_svt_mac l=20n nfin=7 m=4 
MM32 TSMC_26 TSMC_30 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM31 TSMC_22 TSMC_30 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM30 TSMC_30 TSMC_31 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM29 TSMC_31 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM22 TSMC_31 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM9 TSMC_27 TSMC_33 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM8 TSMC_23 TSMC_33 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM7 TSMC_33 TSMC_34 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM5 TSMC_34 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_34 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_25 TSMC_35 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM0 TSMC_24 TSMC_36 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM24 TSMC_21 TSMC_35 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM19 TSMC_20 TSMC_36 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM25 TSMC_35 TSMC_37 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM17 TSMC_36 TSMC_38 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM14 TSMC_37 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM6 TSMC_38 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM15 TSMC_37 TSMC_2 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MP9 TSMC_38 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    PRECHARGE_SB_SD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_PRECHARGE_SB_SD TSMC_1 TSMC_2 TSMC_3 VDDAI VDDI 
MM0_HDM VDDAI TSMC_3 TSMC_1 VDDI pch_svt_mac l=20n nfin=5 m=2 
MP5_HDM TSMC_1 TSMC_3 TSMC_2 VDDI pch_svt_mac l=20n nfin=5 m=1 
MP17_HDM TSMC_2 TSMC_3 VDDAI VDDI pch_svt_mac l=20n nfin=5 m=2 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MCB_2X4_SD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_MCB_2X4_SD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDAI VDDI VSSI TSMC_9 TSMC_10 
XMCB_0<0> TSMC_1 TSMC_5 VDDAI VDDI VSSI TSMC_9 S1ALLSVTSW40W80_BCELL_SD 
XMCB_0<1> TSMC_2 TSMC_6 VDDAI VDDI VSSI TSMC_9 S1ALLSVTSW40W80_BCELL_SD 
XMCB_0<2> TSMC_3 TSMC_7 VDDAI VDDI VSSI TSMC_9 S1ALLSVTSW40W80_BCELL_SD 
XMCB_0<3> TSMC_4 TSMC_8 VDDAI VDDI VSSI TSMC_9 S1ALLSVTSW40W80_BCELL_SD 
XMCB_1<0> TSMC_1 TSMC_5 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW40W80_BCELL_SD 
XMCB_1<1> TSMC_2 TSMC_6 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW40W80_BCELL_SD 
XMCB_1<2> TSMC_3 TSMC_7 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW40W80_BCELL_SD 
XMCB_1<3> TSMC_4 TSMC_8 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW40W80_BCELL_SD 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MIO_M4_SB_BUF
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_MIO_M4_SB_BUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VSSI 
XI8 VSSI VSSI TSMC_6 TSMC_7 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI9 VSSI VSSI TSMC_7 TSMC_4 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI15 VSSI VSSI TSMC_8 TSMC_2 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI14 VSSI VSSI TSMC_9 TSMC_8 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI16 VSSI VSSI TSMC_3 TSMC_6 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI17 VSSI VSSI TSMC_1 TSMC_9 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DIO_TALL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DIO_TALL TSMC_1 TSMC_2 
XDDIO_TALL TSMC_2 TSMC_1 ndio_mac nfin=2 l=2e-07 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    XDRV_STRAP_BT_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_XDRV_STRAP_BT_SB TSMC_1 TSMC_2 VDDI VSSI 
MM0 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=12 m=4 
MM10 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=6 m=12 
MM1 TSMC_2 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=3 m=10 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    RESETD_WTSEL_SB_NEW
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_RESETD_WTSEL_SB_NEW TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ TSMC_3 TSMC_4 
XI87 TSMC_5 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_7 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND5 TSMC_4 TSMC_8 VSSI VSSI VDDHD VDDI TSMC_5 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI84 TSMC_3 TSMC_9 VSSI VSSI VDDHD VDDI TSMC_6 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND0 TSMC_5 TSMC_1 VSSI VSSI VDDHD VDDI TSMC_9 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI89 VSSI VSSI TSMC_7 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI65 VSSI VSSI TSMC_10 TSMC_11 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI83 VSSI VSSI TSMC_11 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI64 VSSI VSSI TSMC_1 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    RESETD_TSEL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_RESETD_TSEL TSMC_1 TSMC_2 TSMC_3 VDDHD VDDI VSSI TSMC_4 
+ TSMC_5 
MM15 TSMC_6 TSMC_1 TSMC_7 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14 TSMC_7 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM25 TSMC_4 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM23 TSMC_4 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM18 TSMC_6 TSMC_1 TSMC_9 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM19 TSMC_9 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM24 TSMC_10 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM21 TSMC_4 TSMC_2 TSMC_10 VSSI nch_svt_mac l=20n nfin=3 m=1 
XI737 VSSI VSSI TSMC_11 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI736 VSSI VSSI TSMC_12 TSMC_11 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND0 TSMC_1 TSMC_5 VSSI VSSI VDDHD VDDI TSMC_8 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI91 TSMC_3 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_12 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    WEBBUF_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_WEBBUF_SB_BASE TSMC_1 TSMC_2 VDDHD VDDI VSSI TSMC_3 
+ TSMC_4 TSMC_5 
MM36 TSMC_6 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM35 TSMC_8 TSMC_2 TSMC_6 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM31 TSMC_9 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=5 m=2 
MM30 TSMC_8 TSMC_3 TSMC_9 VSSI nch_svt_mac l=20n nfin=5 m=1 
MM34 TSMC_10 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM33 TSMC_8 TSMC_1 TSMC_10 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM6 TSMC_8 TSMC_3 TSMC_11 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM32 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
XI25 VSSI VSSI TSMC_8 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI32 VSSI VSSI TSMC_8 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=7 p_l=20n 
XI33 VSSI VSSI TSMC_5 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB4_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 VDDHD VDDI VSSI 
MM15 TSMC_10 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM16 TSMC_10 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM17 TSMC_11 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM18 TSMC_11 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM22 TSMC_11 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM23 TSMC_10 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM24 TSMC_12 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM25 TSMC_13 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_12 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_12 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM2 TSMC_13 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_13 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM19 TSMC_14 TSMC_4 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=2 
MM20 TSMC_10 TSMC_2 TSMC_14 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM21 TSMC_11 TSMC_1 TSMC_14 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM26 TSMC_15 TSMC_5 VSSI VSSI nch_svt_mac l=20n nfin=3 m=4 
MM8 TSMC_16 TSMC_3 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=2 
MM7 TSMC_12 TSMC_2 TSMC_16 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM0 TSMC_13 TSMC_1 TSMC_16 VSSI nch_svt_mac l=20n nfin=3 m=1 
XINV3 VSSI VSSI TSMC_10 TSMC_9 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV2 VSSI VSSI TSMC_11 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV1 VSSI VSSI TSMC_12 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV0 VSSI VSSI TSMC_13 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB1_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VDDHD VDDI VSSI 
MTN1 TSMC_8 TSMC_1 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_9 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MM0 TSMC_8 TSMC_2 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=4 
MM1 TSMC_10 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_8 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=6 
MP5 TSMC_8 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_8 TSMC_1 TSMC_10 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB2_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB2_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD VDDI 
+ VSSI 
MM2 TSMC_6 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_6 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_7 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_7 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM0 TSMC_6 TSMC_1 TSMC_8 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_7 TSMC_2 TSMC_8 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM8 TSMC_8 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=3 m=2 
XINV0 VSSI VSSI TSMC_7 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV1 VSSI VSSI TSMC_6 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_BLEQ_SB_M4
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB1_BLEQ_SB_M4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 VDDHD VDDI VSSI 
MN0 TSMC_1 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=8 m=4 
MTN1 TSMC_7 TSMC_3 TSMC_6 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MM0 TSMC_7 TSMC_4 TSMC_6 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM2 TSMC_2 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=8 m=4 
MP0 TSMC_1 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=6 
MM4 TSMC_7 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM3 TSMC_7 TSMC_3 TSMC_8 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_8 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_2 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=6 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_WLNAD2_SB_X0
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD VDDI VSSI 
MM5 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MTN1 TSMC_9 TSMC_1 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_10 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM0 TSMC_9 TSMC_2 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=6 
MM4 TSMC_8 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MM1 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_9 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=3 
MP5 TSMC_9 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CKBUF_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_CKBUF_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI VSSI 
XINV0 VSSI VSSI TSMC_1 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=7 n_l=20n p_totalM=3 
+ p_nfin=9 p_l=20n 
MM1 TSMC_1 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM34 TSMC_1 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=7 m=2 
MM26 TSMC_5 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=9 m=2 
MM0 TSMC_1 TSMC_4 TSMC_5 VDDI pch_svt_mac l=20n nfin=9 m=2 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    ABUF_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_ABUF_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VSSI 
MM15 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM14 TSMC_3 TSMC_5 TSMC_8 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM9 TSMC_10 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM8 TSMC_3 TSMC_1 TSMC_10 VSSI nch_svt_mac l=20n nfin=4 m=1 
MM13 TSMC_11 TSMC_9 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM12 TSMC_3 TSMC_4 TSMC_11 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM11 TSMC_3 TSMC_1 TSMC_12 TSMC_6 pch_svt_mac l=20n nfin=5 m=1 
MM10 TSMC_12 TSMC_5 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=5 m=2 
XI34 VSSI VSSI TSMC_3 TSMC_9 TSMC_7 TSMC_6 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI35 VSSI VSSI TSMC_3 TSMC_2 TSMC_7 TSMC_6 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    ENBUFB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_ENBUFB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDHD VDDI VSSI 
XI158 TSMC_9 TSMC_9 VSSI VSSI VDDHD VDDI TSMC_10 
+ S1ALLSVTSW40W80_nor2_lvt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM19 TSMC_11 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=6 m=1 
MM2 TSMC_12 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_13 TSMC_8 VDDI VDDI pch_svt_mac l=20n nfin=5 m=1 
MM16 TSMC_13 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=6 m=1 
MM1 TSMC_13 TSMC_2 TSMC_12 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_14 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN200 TSMC_6 TSMC_4 VSSI VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MM4 TSMC_15 TSMC_4 TSMC_14 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_13 TSMC_3 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM20 TSMC_16 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=7 m=1 
MM17 TSMC_13 TSMC_1 TSMC_17 VSSI nch_svt_mac l=20n nfin=4 m=1 
MM18 TSMC_17 TSMC_2 TSMC_16 VSSI nch_svt_mac l=20n nfin=4 m=1 
MN300 TSMC_5 TSMC_4 VSSI VSSI nch_ulvt_mac l=20n nfin=11 m=6 
XI166 VSSI VSSI TSMC_18 TSMC_9 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI148 VSSI VSSI TSMC_4 TSMC_18 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI152 VSSI VSSI TSMC_19 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=4 n_nfin=4 n_l=20n p_totalM=4 
+ p_nfin=8 p_l=20n 
XINV5 VSSI VSSI TSMC_4 TSMC_19 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=3 
+ p_nfin=3 p_l=20n 
XINV4 VSSI VSSI TSMC_10 TSMC_20 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI141 VSSI VSSI TSMC_13 TSMC_4 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=7 n_l=20n p_totalM=3 
+ p_nfin=9 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_WLNAD2_SB_X1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD VDDI VSSI 
MM5 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MTN1 TSMC_9 TSMC_1 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_10 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM0 TSMC_9 TSMC_2 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=6 
MM4 TSMC_8 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MM1 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_9 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=3 
MP5 TSMC_9 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MIO_SB_EDGE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_MIO_SB_EDGE VDDI TSMC_1 TSMC_2 VSSI 
MP0 TSMC_3 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP2 TSMC_4 TSMC_5 VDDI VDDI pch_svt_mac l=20n nfin=3 m=6 
MP7 TSMC_3 TSMC_5 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MN3 VSSI TSMC_3 TSMC_5 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1 VSSI TSMC_3 TSMC_6 VSSI nch_svt_mac l=20n nfin=3 m=5 
MN0 VSSI TSMC_5 TSMC_5 VSSI nch_svt_mac l=20n nfin=3 m=1 
XI18 VSSI VSSI TSMC_4 TSMC_2 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=8 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI393 VSSI VSSI TSMC_6 TSMC_1 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=4 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CKG_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_CKG_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD VDDI 
+ VSSI 
XI58 VSSI VSSI TSMC_6 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM0 TSMC_1 TSMC_7 VDDHD VDDI pch_svt_mac l=16.0n nfin=4 m=1 
MM26 TSMC_1 TSMC_8 VDDHD VDDI pch_svt_mac l=16.0n nfin=4 m=4 
MM1 TSMC_9 TSMC_8 VSSI VSSI nch_svt_mac l=16.0n nfin=8 m=3 
MM34 TSMC_1 TSMC_7 TSMC_9 VSSI nch_svt_mac l=16.0n nfin=8 m=3 
XNAND2 TSMC_2 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_10 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND5 TSMC_4 TSMC_1 VSSI VSSI VDDI VDDI TSMC_7 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND0 TSMC_1 TSMC_5 VSSI VSSI VDDHD VDDI TSMC_11 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND3 TSMC_10 TSMC_11 VSSI VSSI VDDHD VDDI TSMC_6 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND12 TSMC_2 TSMC_3 TSMC_4 VSSI VSSI VDDI VDDI TSMC_8 
+ S1ALLSVTSW40W80_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=10 n_l=16.0n 
+ p_totalM=1 p_nfin=4 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    RESETD_884_M4_SB_NBL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_RESETD_884_M4_SB_NBL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDDHD VDDI VSSI TSMC_12 TSMC_13 
+ TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
XTSEL_WT TSMC_19 TSMC_20 VDDHD VDDI VSSI TSMC_16 TSMC_17 
+ S1ALLSVTSW40W80_RESETD_WTSEL_SB_NEW 
MM10 TSMC_21 TSMC_9 TSMC_11 VDDI pch_svt_mac l=16.0n nfin=3 m=1 
MP0 TSMC_11 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=4 m=3 
MM0 TSMC_22 TSMC_23 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MI537 TSMC_1 TSMC_23 VDDHD VDDI pch_svt_mac l=16.0n nfin=8 m=4 
MM5 TSMC_21 TSMC_24 TSMC_25 VDDI pch_svt_mac l=20n nfin=3 m=1 
XTSEL_READ TSMC_3 TSMC_14 TSMC_15 VDDHD VDDI VSSI TSMC_26 TSMC_27 
+ S1ALLSVTSW40W80_RESETD_TSEL 
MM12 TSMC_21 TSMC_24 TSMC_11 VSSI nch_svt_mac l=16.0n nfin=4 m=2 
MM11 TSMC_1 TSMC_23 VSSI VSSI nch_svt_mac l=16.0n nfin=5 m=4 
MM4 TSMC_21 TSMC_9 TSMC_25 VSSI nch_svt_mac l=20n nfin=4 m=2 
MM1 TSMC_8 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=5 m=1 
XNAND3 TSMC_27 TSMC_26 TSMC_3 VSSI VSSI VDDI VDDI TSMC_23 
+ S1ALLSVTSW40W80_nand3_lvt_mac_pcell_2 n_totalM=2 n_nfin=9 n_l=16.0n 
+ p_totalM=2 p_nfin=3 p_l=16.0n 
XI667 TSMC_19 TSMC_2 TSMC_28 VSSI VSSI VDDHD VDDI TSMC_29 
+ S1ALLSVTSW40W80_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=9 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XI696 TSMC_19 TSMC_20 VSSI VSSI VDDHD VDDI TSMC_30 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI658 TSMC_18 TSMC_1 VSSI VSSI VDDHD VDDI TSMC_31 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI728 TSMC_1 TSMC_32 VSSI VSSI VDDHD VDDI TSMC_25 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI666 TSMC_29 TSMC_33 VSSI VSSI VDDHD VDDI TSMC_34 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XI654 TSMC_31 TSMC_30 VSSI VSSI TSMC_22 VDDI TSMC_8 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI725 VSSI VSSI TSMC_9 TSMC_24 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI730 VSSI VSSI TSMC_35 TSMC_36 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI731 VSSI VSSI TSMC_36 TSMC_37 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI732 VSSI VSSI TSMC_37 TSMC_38 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI733 VSSI VSSI TSMC_38 TSMC_28 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI703 VSSI VSSI TSMC_12 TSMC_35 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI695 VSSI VSSI TSMC_39 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=3 n_nfin=6 n_l=20n p_totalM=4 
+ p_nfin=7 p_l=20n 
XI679 VSSI VSSI TSMC_34 TSMC_40 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=9 n_l=16.0n p_totalM=1 
+ p_nfin=8 p_l=16.0n 
XI693 VSSI VSSI TSMC_3 TSMC_39 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XI713 VSSI VSSI TSMC_21 TSMC_19 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=16.0n p_totalM=2 
+ p_nfin=3 p_l=16.0n 
XI718 VSSI VSSI TSMC_6 TSMC_32 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI686 VSSI VSSI TSMC_41 TSMC_33 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI687 VSSI VSSI TSMC_40 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=8 n_nfin=7 n_l=16.0n p_totalM=8 
+ p_nfin=10 p_l=16.0n 
XI685 VSSI VSSI TSMC_31 TSMC_41 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    COTH_M4_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_COTH_M4_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ VSSI TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
XCKG TSMC_5 TSMC_7 TSMC_8 TSMC_9 TSMC_25 TSMC_16 TSMC_15 VSSI 
+ S1ALLSVTSW40W80_CKG_SB 
XWEBBUF TSMC_3 TSMC_4 TSMC_16 TSMC_15 VSSI TSMC_17 TSMC_18 TSMC_19 
+ S1ALLSVTSW40W80_WEBBUF_SB_BASE 
XRESETD TSMC_1 TSMC_2 TSMC_5 TSMC_6 TSMC_26 TSMC_7 TSMC_21 TSMC_25 TSMC_12 
+ TSMC_13 TSMC_14 TSMC_16 TSMC_15 VSSI TSMC_19 TSMC_20 TSMC_10 TSMC_11 
+ TSMC_22 TSMC_23 TSMC_24 S1ALLSVTSW40W80_RESETD_884_M4_SB_NBL 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_Y_M4_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB1_Y_M4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VDDHD VDDI VSSI 
MM6 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=9 m=9 
MTN1 TSMC_9 TSMC_1 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_10 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM0 TSMC_9 TSMC_2 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM7 TSMC_8 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=7 m=6 
MM3 TSMC_9 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP5 TSMC_9 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM1 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM2 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_DCLK_M4_SB_V2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DECB1_DCLK_M4_SB_V2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD VDDI VSSI 
MM2 TSMC_4 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=5 
MTN1 TSMC_8 TSMC_1 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_9 TSMC_7 TSMC_6 VSSI nch_ulvt_mac l=20n nfin=6 m=4 
MM0 TSMC_8 TSMC_2 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=6 m=4 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=5 
MM4 TSMC_4 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=8 
MM1 TSMC_10 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_8 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=8 
MP5 TSMC_8 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM5 TSMC_8 TSMC_1 TSMC_10 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CDEC_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_CDEC_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 VSSI TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 
XPREDEC_Y<0> TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_47 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_45 TSMC_44 VSSI S1ALLSVTSW40W80_DECB4_SB 
XPREDEC_Y<1> TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_48 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_45 TSMC_44 VSSI S1ALLSVTSW40W80_DECB4_SB 
XIPDEC_X1<0> TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 
+ TSMC_83 TSMC_45 TSMC_44 VSSI S1ALLSVTSW40W80_DECB4_SB 
XIPDEC_X1<1> TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_45 TSMC_44 VSSI S1ALLSVTSW40W80_DECB4_SB 
XIPDEC_X0<0> TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_45 TSMC_44 VSSI S1ALLSVTSW40W80_DECB4_SB 
XIPDEC_X0<1> TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_45 TSMC_44 VSSI S1ALLSVTSW40W80_DECB4_SB 
XIDEC_X2<0> TSMC_8 TSMC_10 TSMC_28 TSMC_40 TSMC_103 TSMC_41 TSMC_104 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_SB 
XIDEC_X2<1> TSMC_8 TSMC_10 TSMC_29 TSMC_40 TSMC_103 TSMC_41 TSMC_105 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_SB 
XIDEC_X2<2> TSMC_8 TSMC_10 TSMC_30 TSMC_40 TSMC_103 TSMC_41 TSMC_106 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_SB 
XIDEC_X2<3> TSMC_8 TSMC_10 TSMC_31 TSMC_40 TSMC_103 TSMC_41 TSMC_107 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_SB 
XI381<0> TSMC_108 TSMC_109 TSMC_110 TSMC_104 TSMC_105 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW40W80_DECB2_SB 
XI381<1> TSMC_108 TSMC_109 TSMC_111 TSMC_106 TSMC_107 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW40W80_DECB2_SB 
XDECB1_BLEQ TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_112 TSMC_113 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW40W80_DECB1_BLEQ_SB_M4 
XIDEC_X0<0> TSMC_9 TSMC_10 TSMC_12 TSMC_112 TSMC_113 TSMC_41 TSMC_94 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XIDEC_X0<1> TSMC_9 TSMC_10 TSMC_13 TSMC_112 TSMC_113 TSMC_41 TSMC_95 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XIDEC_X0<2> TSMC_9 TSMC_10 TSMC_14 TSMC_112 TSMC_113 TSMC_41 TSMC_96 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XIDEC_X0<3> TSMC_9 TSMC_10 TSMC_15 TSMC_112 TSMC_113 TSMC_41 TSMC_97 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XIDEC_X0<4> TSMC_9 TSMC_10 TSMC_16 TSMC_112 TSMC_113 TSMC_41 TSMC_99 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XIDEC_X0<5> TSMC_9 TSMC_10 TSMC_17 TSMC_112 TSMC_113 TSMC_41 TSMC_100 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XIDEC_X0<6> TSMC_9 TSMC_10 TSMC_18 TSMC_112 TSMC_113 TSMC_41 TSMC_101 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XIDEC_X0<7> TSMC_9 TSMC_10 TSMC_19 TSMC_112 TSMC_113 TSMC_41 TSMC_102 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X0 
XCKBUF TSMC_4 TSMC_5 TSMC_9 TSMC_11 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW40W80_CKBUF_SB 
XABUF_Y<0> TSMC_57 TSMC_63 TSMC_64 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_Y<1> TSMC_58 TSMC_65 TSMC_66 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<3> TSMC_52 TSMC_75 TSMC_76 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<4> TSMC_53 TSMC_77 TSMC_78 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<5> TSMC_54 TSMC_79 TSMC_84 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<6> TSMC_55 TSMC_108 TSMC_109 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<7> TSMC_56 TSMC_110 TSMC_111 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<0> TSMC_49 TSMC_89 TSMC_90 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<1> TSMC_50 TSMC_91 TSMC_92 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XABUF_X<2> TSMC_51 TSMC_93 TSMC_98 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW40W80_ABUF_SB_BASE 
XIDEC_Y<0> TSMC_9 TSMC_10 TSMC_32 TSMC_112 TSMC_113 TSMC_41 TSMC_67 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_Y<1> TSMC_9 TSMC_10 TSMC_33 TSMC_112 TSMC_113 TSMC_41 TSMC_68 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_Y<2> TSMC_9 TSMC_10 TSMC_34 TSMC_112 TSMC_113 TSMC_41 TSMC_69 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_Y<3> TSMC_9 TSMC_10 TSMC_35 TSMC_112 TSMC_113 TSMC_41 TSMC_70 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_Y<4> TSMC_9 TSMC_11 TSMC_36 TSMC_112 TSMC_113 TSMC_41 TSMC_71 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_Y<5> TSMC_9 TSMC_11 TSMC_37 TSMC_112 TSMC_113 TSMC_41 TSMC_72 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_Y<6> TSMC_9 TSMC_11 TSMC_38 TSMC_112 TSMC_113 TSMC_41 TSMC_73 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_Y<7> TSMC_9 TSMC_11 TSMC_39 TSMC_112 TSMC_113 TSMC_41 TSMC_74 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_Y_M4_SB 
XIDEC_CKD TSMC_9 TSMC_10 TSMC_6 TSMC_7 TSMC_112 TSMC_113 TSMC_48 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_DCLK_M4_SB_V2 
XIDEC_X1<0> TSMC_9 TSMC_10 TSMC_20 TSMC_112 TSMC_113 TSMC_41 TSMC_80 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XIDEC_X1<1> TSMC_9 TSMC_10 TSMC_21 TSMC_112 TSMC_113 TSMC_41 TSMC_81 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XIDEC_X1<2> TSMC_9 TSMC_10 TSMC_22 TSMC_112 TSMC_113 TSMC_41 TSMC_82 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XIDEC_X1<3> TSMC_9 TSMC_10 TSMC_23 TSMC_112 TSMC_113 TSMC_41 TSMC_83 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XIDEC_X1<4> TSMC_9 TSMC_10 TSMC_24 TSMC_112 TSMC_113 TSMC_41 TSMC_85 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XIDEC_X1<5> TSMC_9 TSMC_10 TSMC_25 TSMC_112 TSMC_113 TSMC_41 TSMC_86 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XIDEC_X1<6> TSMC_9 TSMC_10 TSMC_26 TSMC_112 TSMC_113 TSMC_41 TSMC_87 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XIDEC_X1<7> TSMC_9 TSMC_10 TSMC_27 TSMC_112 TSMC_113 TSMC_41 TSMC_88 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_DECB1_WLNAD2_SB_X1 
XCEBBUF TSMC_3 TSMC_4 TSMC_5 TSMC_40 TSMC_113 TSMC_103 TSMC_112 TSMC_43 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW40W80_ENBUFB_BASE 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CNT_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_CNT_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 VSSI TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 
XCOTHERS TSMC_3 TSMC_3 TSMC_65 TSMC_66 TSMC_7 TSMC_67 TSMC_8 TSMC_68 TSMC_69 
+ TSMC_42 TSMC_43 TSMC_45 TSMC_70 TSMC_46 TSMC_47 TSMC_47 VSSI TSMC_48 
+ TSMC_71 TSMC_49 TSMC_44 TSMC_72 TSMC_50 TSMC_51 TSMC_52 
+ S1ALLSVTSW40W80_COTH_M4_BASE 
Xcdec TSMC_1 TSMC_2 TSMC_4 TSMC_65 TSMC_66 TSMC_5 TSMC_6 TSMC_7 TSMC_67 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_68 TSMC_73 TSMC_74 
+ TSMC_69 TSMC_47 TSMC_47 VSSI TSMC_75 TSMC_71 TSMC_49 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_76 TSMC_77 S1ALLSVTSW40W80_CDEC_M4_SB_BASE 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DIN_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DIN_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI 
+ VSSI TSMC_5 TSMC_6 
MM6 TSMC_7 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM4 TSMC_9 TSMC_10 TSMC_11 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM35 TSMC_12 TSMC_13 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM41 TSMC_14 TSMC_13 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN33 TSMC_7 TSMC_15 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM19 TSMC_16 TSMC_1 TSMC_17 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM1 VSSI TSMC_8 TSMC_18 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM12 TSMC_16 TSMC_10 TSMC_14 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM5 VSSI TSMC_19 TSMC_11 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM9 TSMC_20 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM42 TSMC_17 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM34 TSMC_9 TSMC_3 TSMC_18 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM8 TSMC_20 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM39 TSMC_22 TSMC_10 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM26 VDDHD TSMC_10 TSMC_23 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_24 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MM2 VDDHD TSMC_19 TSMC_25 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM33 TSMC_21 TSMC_13 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM36 TSMC_15 TSMC_13 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_9 TSMC_8 TSMC_25 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM14 TSMC_20 TSMC_21 TSMC_24 VDDI pch_svt_mac l=20n nfin=3 m=2 
MM0 TSMC_9 TSMC_3 TSMC_23 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM51 TSMC_7 TSMC_15 TSMC_24 VDDI pch_svt_mac l=20n nfin=3 m=2 
MM16 TSMC_16 TSMC_8 TSMC_26 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM15 TSMC_16 TSMC_1 TSMC_22 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM40 TSMC_26 TSMC_13 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
XI395 TSMC_12 VSSI TSMC_9 TSMC_21 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI295 TSMC_4 VSSI TSMC_7 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=3 n_nfin=9 n_l=20n p_totalM=3 
+ p_nfin=2 p_l=20n 
XI341 VSSI VSSI TSMC_2 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI396 TSMC_12 VSSI TSMC_19 TSMC_15 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI277 VSSI VSSI TSMC_16 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI339 TSMC_4 VSSI TSMC_20 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=3 n_nfin=9 n_l=20n p_totalM=3 
+ p_nfin=2 p_l=20n 
XI386 VSSI VSSI TSMC_8 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XINV04 VSSI VSSI TSMC_9 TSMC_19 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DOUT_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DOUT_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD VDDI 
+ VSSI 
MP11 TSMC_6 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM12 TSMC_6 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM9 TSMC_8 TSMC_7 TSMC_6 VDDI pch_svt_mac l=20n nfin=5 m=2 
MM17 TSMC_9 TSMC_10 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM8 TSMC_8 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MP14 TSMC_6 TSMC_12 TSMC_3 VDDI pch_svt_mac l=20n nfin=5 m=1 
MP13 TSMC_8 TSMC_12 TSMC_2 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM14_SA TSMC_13 TSMC_8 VDDHD VDDI pch_lvt_mac l=20n nfin=6 m=1 
MP2 TSMC_8 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MP10 TSMC_4 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=4 m=4 
MM35_SA TSMC_14 TSMC_6 VDDHD VDDI pch_lvt_mac l=20n nfin=6 m=1 
MM24_SA TSMC_15 TSMC_16 TSMC_14 VDDI pch_lvt_mac l=20n nfin=6 m=1 
MM20 TSMC_11 TSMC_17 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM23_SA TSMC_9 TSMC_16 TSMC_13 VDDI pch_lvt_mac l=20n nfin=6 m=1 
MM31_SA TSMC_18 TSMC_6 VSSI VSSI nch_lvt_mac l=20n nfin=3 m=1 
MN1 TSMC_6 TSMC_8 TSMC_19 VSSI nch_svt_mac l=20n nfin=10 m=4 
MM7 TSMC_19 TSMC_10 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM6 TSMC_8 TSMC_6 TSMC_19 VSSI nch_svt_mac l=20n nfin=10 m=4 
MM15_SA TSMC_20 TSMC_8 VSSI VSSI nch_lvt_mac l=20n nfin=3 m=1 
MM13_SA TSMC_9 TSMC_10 TSMC_20 VSSI nch_lvt_mac l=20n nfin=3 m=1 
MM18 TSMC_9 TSMC_16 TSMC_21 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN5 TSMC_4 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=4 m=4 
MM29_SA TSMC_15 TSMC_10 TSMC_18 VSSI nch_lvt_mac l=20n nfin=3 m=1 
MM21 TSMC_21 TSMC_17 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
XIPGB0 TSMC_22 TSMC_16 TSMC_7 VSSI VSSI VDDHD VDDI TSMC_12 
+ S1ALLSVTSW40W80_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI159 TSMC_16 TSMC_23 VSSI VSSI VDDHD VDDI TSMC_7 
+ S1ALLSVTSW40W80_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI185 VSSI VSSI TSMC_16 TSMC_24 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI203 VSSI VSSI TSMC_25 TSMC_23 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI184 VSSI VSSI TSMC_10 TSMC_16 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI161 VSSI VSSI TSMC_26 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI194 VSSI VSSI TSMC_5 TSMC_26 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI186 VSSI VSSI TSMC_24 TSMC_22 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI201 VSSI VSSI TSMC_1 TSMC_25 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI163 VSSI VSSI TSMC_9 TSMC_17 VDDHD VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    YPASS_M4_SB_NBL_V2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_YPASS_M4_SB_NBL_V2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 VDDI VSSI TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
XI250<4> TSMC_13 VSSI TSMC_20 TSMC_24 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI250<5> TSMC_13 VSSI TSMC_21 TSMC_25 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI250<6> TSMC_13 VSSI TSMC_22 TSMC_26 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI250<7> TSMC_13 VSSI TSMC_23 TSMC_27 VDDI VDDI 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MN18<0> TSMC_5 TSMC_24 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN18<1> TSMC_6 TSMC_25 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN18<2> TSMC_7 TSMC_26 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN18<3> TSMC_8 TSMC_27 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<0> TSMC_1 TSMC_24 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<1> TSMC_2 TSMC_25 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<2> TSMC_3 TSMC_26 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<3> TSMC_4 TSMC_27 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MM4 TSMC_10 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM0 TSMC_28 TSMC_10 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM5 TSMC_10 TSMC_9 VDDI VDDI pch_svt_mac l=20n nfin=4 m=1 
MP10<0> TSMC_12 TSMC_16 TSMC_5 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP10<1> TSMC_12 TSMC_17 TSMC_6 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP10<2> TSMC_12 TSMC_18 TSMC_7 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP10<3> TSMC_12 TSMC_19 TSMC_8 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP3_HDM TSMC_12 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP22_HDM VDDI TSMC_28 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<0> TSMC_11 TSMC_16 TSMC_1 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<1> TSMC_11 TSMC_17 TSMC_2 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<2> TSMC_11 TSMC_18 TSMC_3 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<3> TSMC_11 TSMC_19 TSMC_4 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_28 TSMC_10 VDDI VDDI pch_svt_mac l=20n nfin=4 m=3 
MM14<0> TSMC_1 TSMC_5 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14<1> TSMC_2 TSMC_6 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14<2> TSMC_3 TSMC_7 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14<3> TSMC_4 TSMC_8 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<0> TSMC_5 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<1> TSMC_6 TSMC_2 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<2> TSMC_7 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<3> TSMC_8 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
XPRECHARGE<0> TSMC_1 TSMC_5 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW40W80_PRECHARGE_SB_SD 
XPRECHARGE<1> TSMC_2 TSMC_6 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW40W80_PRECHARGE_SB_SD 
XPRECHARGE<2> TSMC_3 TSMC_7 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW40W80_PRECHARGE_SB_SD 
XPRECHARGE<3> TSMC_4 TSMC_8 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW40W80_PRECHARGE_SB_SD 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MIO_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_MIO_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 VSSI TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
XDIN TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_16 TSMC_16 VSSI TSMC_25 TSMC_26 
+ S1ALLSVTSW40W80_DIN_M4_SB_BASE 
XDOUT TSMC_27 TSMC_28 TSMC_29 TSMC_14 TSMC_15 TSMC_16 TSMC_16 VSSI 
+ S1ALLSVTSW40W80_DOUT_SB 
XYPASS TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_27 
+ TSMC_28 TSMC_29 TSMC_13 TSMC_16 VSSI TSMC_25 TSMC_26 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ S1ALLSVTSW40W80_YPASS_M4_SB_NBL_V2 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CNT_M4_SB_BUF
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_CNT_M4_SB_BUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VSSI 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
XI32 VSSI VSSI TSMC_32 TSMC_4 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=10 n_l=20n p_totalM=2 
+ p_nfin=10 p_l=20n 
XI31 VSSI VSSI TSMC_3 TSMC_32 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=10 n_l=20n p_totalM=1 
+ p_nfin=10 p_l=20n 
XWEB_INV VSSI VSSI TSMC_6 TSMC_7 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI29<0> VSSI VSSI TSMC_24 TSMC_28 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI29<1> VSSI VSSI TSMC_25 TSMC_29 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI30 VSSI VSSI TSMC_1 TSMC_2 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
XI28<0> VSSI VSSI TSMC_8 TSMC_16 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<1> VSSI VSSI TSMC_9 TSMC_17 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<2> VSSI VSSI TSMC_10 TSMC_18 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<3> VSSI VSSI TSMC_11 TSMC_19 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<4> VSSI VSSI TSMC_12 TSMC_20 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<5> VSSI VSSI TSMC_13 TSMC_21 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<6> VSSI VSSI TSMC_14 TSMC_22 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<7> VSSI VSSI TSMC_15 TSMC_23 TSMC_5 TSMC_5 
+ S1ALLSVTSW40W80_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DIODE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_DIODE TSMC_1 TSMC_2 TSMC_3 
MMDIODE TSMC_1 TSMC_2 TSMC_1 TSMC_3 nch_lvt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    LOGIC_D0907_TRKWL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_LOGIC_D0907_TRKWL TSMC_1 TSMC_2 
MM2 TSMC_1 TSMC_2 TSMC_1 TSMC_1 nch_svt_mac l=20n nfin=4 m=1 
MM1 TSMC_1 TSMC_2 TSMC_1 TSMC_1 nch_svt_mac l=20n nfin=4 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MCB_D0907_ONCELL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW40W80_MCB_D0907_ONCELL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
Mpd11 TSMC_9 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg21 TSMC_11 TSMC_7 TSMC_10 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_12 TSMC_13 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg11 TSMC_1 TSMC_2 TSMC_9 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_13 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_13 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_11 TSMC_8 TSMC_12 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpu11 TSMC_9 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_13 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS




**** End of leaf cells

.SUBCKT S1ALLSVTSW40W80_MCB_ARR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDAI VDDI VSSI TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 
XMCB_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_9 TSMC_10 S1ALLSVTSW40W80_MCB_2X4_SD 
XMCB_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_11 TSMC_12 S1ALLSVTSW40W80_MCB_2X4_SD 
XMCB_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_13 TSMC_14 S1ALLSVTSW40W80_MCB_2X4_SD 
XMCB_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_15 TSMC_16 S1ALLSVTSW40W80_MCB_2X4_SD 
XMCB_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_17 TSMC_18 S1ALLSVTSW40W80_MCB_2X4_SD 
XMCB_5 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_19 TSMC_20 S1ALLSVTSW40W80_MCB_2X4_SD 
XMCB_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_21 TSMC_22 S1ALLSVTSW40W80_MCB_2X4_SD 
XMCB_7 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_2X4_SD 
.ENDS

.SUBCKT S1ALLSVTSW40W80_TRACKING_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 VDDI VSSI TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 
XTKBL_ON_CELL_0 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_273 
+ TSMC_274 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_1 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_271 
+ TSMC_272 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_2 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_269 
+ TSMC_270 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_3 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_267 
+ TSMC_268 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_4 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_265 
+ TSMC_266 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_5 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_263 
+ TSMC_264 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_6 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_261 
+ TSMC_262 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_7 TSMC_257 TSMC_275 TSMC_275 VDDI TSMC_258 VSSI TSMC_259 
+ TSMC_260 S1ALLSVTSW40W80_MCB_D0907_ONCELL 
XTRKWL_CELL_0 VSSI TSMC_275 S1ALLSVTSW40W80_LOGIC_D0907_TRKWL 
XTRKWL_CELL_1 VSSI TSMC_275 S1ALLSVTSW40W80_LOGIC_D0907_TRKWL 
XTRKWL_CELL_2 VSSI TSMC_275 S1ALLSVTSW40W80_LOGIC_D0907_TRKWL 
.ENDS

.SUBCKT S1ALLSVTSW40W80_MIO_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 VSSI TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
XMIO_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_24 TSMC_11 TSMC_25 VSSI TSMC_13 TSMC_14 TSMC_15 VSSI TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ S1ALLSVTSW40W80_MIO_M4_SB_BASE 
XMIO_MX_SB_BUF TSMC_10 TSMC_24 TSMC_12 TSMC_25 TSMC_15 VSSI 
+ S1ALLSVTSW40W80_MIO_M4_SB_BUF 
.ENDS

.SUBCKT S1ALLSVTSW40W80_CNT_M4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 VSSI TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
XCNT_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_62 TSMC_5 TSMC_6 TSMC_63 TSMC_7 
+ TSMC_64 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 VSSI TSMC_65 
+ TSMC_66 TSMC_47 TSMC_48 TSMC_49 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ S1ALLSVTSW40W80_CNT_M4_SB_BASE 
XCNT_MX_SB_BUF TSMC_4 TSMC_62 TSMC_7 TSMC_64 TSMC_45 VSSI TSMC_46 TSMC_65 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_58 
+ TSMC_59 TSMC_60 TSMC_61 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ S1ALLSVTSW40W80_CNT_M4_SB_BUF 
.ENDS

.SUBCKT TS1N16FFCLLSVTA64X128M4SW D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] D[8] 
+ D[9] D[10] D[11] D[12] D[13] D[14] D[15] D[16] D[17] D[18] D[19] D[20] D[21] 
+ D[22] D[23] D[24] D[25] D[26] D[27] D[28] D[29] D[30] D[31] D[32] D[33] D[34] 
+ D[35] D[36] D[37] D[38] D[39] D[40] D[41] D[42] D[43] D[44] D[45] D[46] D[47] 
+ D[48] D[49] D[50] D[51] D[52] D[53] D[54] D[55] D[56] D[57] D[58] D[59] D[60] 
+ D[61] D[62] D[63] D[64] D[65] D[66] D[67] D[68] D[69] D[70] D[71] D[72] D[73] 
+ D[74] D[75] D[76] D[77] D[78] D[79] D[80] D[81] D[82] D[83] D[84] D[85] D[86] 
+ D[87] D[88] D[89] D[90] D[91] D[92] D[93] D[94] D[95] D[96] D[97] D[98] D[99] 
+ D[100] D[101] D[102] D[103] D[104] D[105] D[106] D[107] D[108] D[109] D[110] 
+ D[111] D[112] D[113] D[114] D[115] D[116] D[117] D[118] D[119] D[120] D[121] 
+ D[122] D[123] D[124] D[125] D[126] D[127] BWEB[0] BWEB[1] BWEB[2] BWEB[3] 
+ BWEB[4] BWEB[5] BWEB[6] BWEB[7] BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12] 
+ BWEB[13] BWEB[14] BWEB[15] BWEB[16] BWEB[17] BWEB[18] BWEB[19] BWEB[20] 
+ BWEB[21] BWEB[22] BWEB[23] BWEB[24] BWEB[25] BWEB[26] BWEB[27] BWEB[28] 
+ BWEB[29] BWEB[30] BWEB[31] BWEB[32] BWEB[33] BWEB[34] BWEB[35] BWEB[36] 
+ BWEB[37] BWEB[38] BWEB[39] BWEB[40] BWEB[41] BWEB[42] BWEB[43] BWEB[44] 
+ BWEB[45] BWEB[46] BWEB[47] BWEB[48] BWEB[49] BWEB[50] BWEB[51] BWEB[52] 
+ BWEB[53] BWEB[54] BWEB[55] BWEB[56] BWEB[57] BWEB[58] BWEB[59] BWEB[60] 
+ BWEB[61] BWEB[62] BWEB[63] BWEB[64] BWEB[65] BWEB[66] BWEB[67] BWEB[68] 
+ BWEB[69] BWEB[70] BWEB[71] BWEB[72] BWEB[73] BWEB[74] BWEB[75] BWEB[76] 
+ BWEB[77] BWEB[78] BWEB[79] BWEB[80] BWEB[81] BWEB[82] BWEB[83] BWEB[84] 
+ BWEB[85] BWEB[86] BWEB[87] BWEB[88] BWEB[89] BWEB[90] BWEB[91] BWEB[92] 
+ BWEB[93] BWEB[94] BWEB[95] BWEB[96] BWEB[97] BWEB[98] BWEB[99] BWEB[100] 
+ BWEB[101] BWEB[102] BWEB[103] BWEB[104] BWEB[105] BWEB[106] BWEB[107] 
+ BWEB[108] BWEB[109] BWEB[110] BWEB[111] BWEB[112] BWEB[113] BWEB[114] 
+ BWEB[115] BWEB[116] BWEB[117] BWEB[118] BWEB[119] BWEB[120] BWEB[121] 
+ BWEB[122] BWEB[123] BWEB[124] BWEB[125] BWEB[126] BWEB[127] A[0] A[1] A[2] 
+ A[3] A[4] A[5] Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] Q[11] 
+ Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18] Q[19] Q[20] Q[21] Q[22] Q[23] Q[24] 
+ Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] Q[32] Q[33] Q[34] Q[35] Q[36] Q[37] 
+ Q[38] Q[39] Q[40] Q[41] Q[42] Q[43] Q[44] Q[45] Q[46] Q[47] Q[48] Q[49] Q[50] 
+ Q[51] Q[52] Q[53] Q[54] Q[55] Q[56] Q[57] Q[58] Q[59] Q[60] Q[61] Q[62] Q[63] 
+ Q[64] Q[65] Q[66] Q[67] Q[68] Q[69] Q[70] Q[71] Q[72] Q[73] Q[74] Q[75] Q[76] 
+ Q[77] Q[78] Q[79] Q[80] Q[81] Q[82] Q[83] Q[84] Q[85] Q[86] Q[87] Q[88] Q[89] 
+ Q[90] Q[91] Q[92] Q[93] Q[94] Q[95] Q[96] Q[97] Q[98] Q[99] Q[100] Q[101] 
+ Q[102] Q[103] Q[104] Q[105] Q[106] Q[107] Q[108] Q[109] Q[110] Q[111] Q[112] 
+ Q[113] Q[114] Q[115] Q[116] Q[117] Q[118] Q[119] Q[120] Q[121] Q[122] Q[123] 
+ Q[124] Q[125] Q[126] Q[127] CEB CLK WEB RTSEL[1] RTSEL[0] WTSEL[1] WTSEL[0] 
+ VDD VSS 
XMCB16X4_L_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDD VDD 
+ VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_1 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_2 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_3 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_4 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_5 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_6 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_7 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_8 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_9 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_10 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 
+ TSMC_104 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_11 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_12 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 
+ TSMC_120 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_13 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 
+ TSMC_128 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_14 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 
+ TSMC_136 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_15 TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 
+ TSMC_144 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_16 TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_17 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_18 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 
+ TSMC_168 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_19 TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 
+ TSMC_176 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_20 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_21 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 
+ TSMC_192 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_22 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 
+ TSMC_200 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_23 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_24 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_25 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_26 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 
+ TSMC_231 TSMC_232 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_27 TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 
+ TSMC_239 TSMC_240 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_28 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_247 TSMC_248 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_29 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 
+ TSMC_255 TSMC_256 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_30 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 
+ TSMC_263 TSMC_264 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_31 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 
+ TSMC_271 TSMC_272 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_32 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 
+ TSMC_279 TSMC_280 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_33 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 
+ TSMC_287 TSMC_288 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_34 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 
+ TSMC_295 TSMC_296 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_35 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 
+ TSMC_303 TSMC_304 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_36 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 
+ TSMC_311 TSMC_312 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_37 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 
+ TSMC_319 TSMC_320 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_38 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 
+ TSMC_327 TSMC_328 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_39 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 
+ TSMC_335 TSMC_336 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_40 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 
+ TSMC_343 TSMC_344 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_41 TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 
+ TSMC_351 TSMC_352 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_42 TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 
+ TSMC_359 TSMC_360 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_43 TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 
+ TSMC_367 TSMC_368 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_44 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 
+ TSMC_375 TSMC_376 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_45 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_46 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 
+ TSMC_391 TSMC_392 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_47 TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 
+ TSMC_399 TSMC_400 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_48 TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_407 TSMC_408 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_49 TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 
+ TSMC_415 TSMC_416 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_50 TSMC_417 TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 
+ TSMC_423 TSMC_424 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_51 TSMC_425 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 
+ TSMC_431 TSMC_432 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_52 TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 
+ TSMC_439 TSMC_440 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_53 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 
+ TSMC_447 TSMC_448 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_54 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_55 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 
+ TSMC_463 TSMC_464 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_56 TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 
+ TSMC_471 TSMC_472 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_57 TSMC_473 TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 
+ TSMC_479 TSMC_480 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_58 TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 
+ TSMC_487 TSMC_488 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_59 TSMC_489 TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 
+ TSMC_495 TSMC_496 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_60 TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 
+ TSMC_503 TSMC_504 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_61 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_62 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 
+ TSMC_519 TSMC_520 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_L_63 TSMC_521 TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 
+ TSMC_527 TSMC_528 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_64 TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 
+ TSMC_535 TSMC_536 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_65 TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 
+ TSMC_559 TSMC_560 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_66 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_67 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 TSMC_576 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_68 TSMC_577 TSMC_578 TSMC_579 TSMC_580 TSMC_581 TSMC_582 
+ TSMC_583 TSMC_584 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_69 TSMC_585 TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 
+ TSMC_591 TSMC_592 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_70 TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_71 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 
+ TSMC_607 TSMC_608 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_72 TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 
+ TSMC_615 TSMC_616 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_73 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_74 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_75 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 
+ TSMC_639 TSMC_640 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_76 TSMC_641 TSMC_642 TSMC_643 TSMC_644 TSMC_645 TSMC_646 
+ TSMC_647 TSMC_648 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_77 TSMC_649 TSMC_650 TSMC_651 TSMC_652 TSMC_653 TSMC_654 
+ TSMC_655 TSMC_656 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_78 TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 
+ TSMC_663 TSMC_664 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_79 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 
+ TSMC_671 TSMC_672 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_80 TSMC_673 TSMC_674 TSMC_675 TSMC_676 TSMC_677 TSMC_678 
+ TSMC_679 TSMC_680 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_81 TSMC_681 TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 
+ TSMC_687 TSMC_688 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_82 TSMC_689 TSMC_690 TSMC_691 TSMC_692 TSMC_693 TSMC_694 
+ TSMC_695 TSMC_696 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_83 TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_701 TSMC_702 
+ TSMC_703 TSMC_704 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_84 TSMC_705 TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 
+ TSMC_711 TSMC_712 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_85 TSMC_713 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 
+ TSMC_719 TSMC_720 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_86 TSMC_721 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_727 TSMC_728 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_87 TSMC_729 TSMC_730 TSMC_731 TSMC_732 TSMC_733 TSMC_734 
+ TSMC_735 TSMC_736 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_88 TSMC_737 TSMC_738 TSMC_739 TSMC_740 TSMC_741 TSMC_742 
+ TSMC_743 TSMC_744 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_89 TSMC_745 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 
+ TSMC_751 TSMC_752 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_90 TSMC_753 TSMC_754 TSMC_755 TSMC_756 TSMC_757 TSMC_758 
+ TSMC_759 TSMC_760 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_91 TSMC_761 TSMC_762 TSMC_763 TSMC_764 TSMC_765 TSMC_766 
+ TSMC_767 TSMC_768 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_92 TSMC_769 TSMC_770 TSMC_771 TSMC_772 TSMC_773 TSMC_774 
+ TSMC_775 TSMC_776 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_93 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_782 
+ TSMC_783 TSMC_784 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_94 TSMC_785 TSMC_786 TSMC_787 TSMC_788 TSMC_789 TSMC_790 
+ TSMC_791 TSMC_792 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_95 TSMC_793 TSMC_794 TSMC_795 TSMC_796 TSMC_797 TSMC_798 
+ TSMC_799 TSMC_800 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_96 TSMC_801 TSMC_802 TSMC_803 TSMC_804 TSMC_805 TSMC_806 
+ TSMC_807 TSMC_808 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_97 TSMC_809 TSMC_810 TSMC_811 TSMC_812 TSMC_813 TSMC_814 
+ TSMC_815 TSMC_816 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_98 TSMC_817 TSMC_818 TSMC_819 TSMC_820 TSMC_821 TSMC_822 
+ TSMC_823 TSMC_824 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_99 TSMC_825 TSMC_826 TSMC_827 TSMC_828 TSMC_829 TSMC_830 
+ TSMC_831 TSMC_832 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_100 TSMC_833 TSMC_834 TSMC_835 TSMC_836 TSMC_837 TSMC_838 
+ TSMC_839 TSMC_840 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_101 TSMC_841 TSMC_842 TSMC_843 TSMC_844 TSMC_845 TSMC_846 
+ TSMC_847 TSMC_848 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_102 TSMC_849 TSMC_850 TSMC_851 TSMC_852 TSMC_853 TSMC_854 
+ TSMC_855 TSMC_856 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_103 TSMC_857 TSMC_858 TSMC_859 TSMC_860 TSMC_861 TSMC_862 
+ TSMC_863 TSMC_864 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_104 TSMC_865 TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 
+ TSMC_871 TSMC_872 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_105 TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 
+ TSMC_879 TSMC_880 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_106 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 
+ TSMC_887 TSMC_888 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_107 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_108 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 TSMC_902 
+ TSMC_903 TSMC_904 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_109 TSMC_905 TSMC_906 TSMC_907 TSMC_908 TSMC_909 TSMC_910 
+ TSMC_911 TSMC_912 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_110 TSMC_913 TSMC_914 TSMC_915 TSMC_916 TSMC_917 TSMC_918 
+ TSMC_919 TSMC_920 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_111 TSMC_921 TSMC_922 TSMC_923 TSMC_924 TSMC_925 TSMC_926 
+ TSMC_927 TSMC_928 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_112 TSMC_929 TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 
+ TSMC_935 TSMC_936 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_113 TSMC_937 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 
+ TSMC_943 TSMC_944 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_114 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_115 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 TSMC_958 
+ TSMC_959 TSMC_960 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_116 TSMC_961 TSMC_962 TSMC_963 TSMC_964 TSMC_965 TSMC_966 
+ TSMC_967 TSMC_968 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_117 TSMC_969 TSMC_970 TSMC_971 TSMC_972 TSMC_973 TSMC_974 
+ TSMC_975 TSMC_976 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_118 TSMC_977 TSMC_978 TSMC_979 TSMC_980 TSMC_981 TSMC_982 
+ TSMC_983 TSMC_984 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_119 TSMC_985 TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 
+ TSMC_991 TSMC_992 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_120 TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 
+ TSMC_999 TSMC_1000 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_121 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_122 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 TSMC_1013 TSMC_1014 
+ TSMC_1015 TSMC_1016 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_123 TSMC_1017 TSMC_1018 TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 
+ TSMC_1023 TSMC_1024 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_124 TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_125 TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 TSMC_1037 TSMC_1038 
+ TSMC_1039 TSMC_1040 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_126 TSMC_1041 TSMC_1042 TSMC_1043 TSMC_1044 TSMC_1045 TSMC_1046 
+ TSMC_1047 TSMC_1048 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XMCB16X4_R_127 TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 
+ TSMC_1055 TSMC_1056 VDD VDD VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ S1ALLSVTSW40W80_MCB_ARR 
XXDRV_STRAP_BT_SB_0 TSMC_1057 TSMC_1058 VDD VSS 
+ S1ALLSVTSW40W80_XDRV_STRAP_BT_SB 
XXDRV_LA512_SB_0 TSMC_1059 TSMC_1060 TSMC_1061 TSMC_1062 TSMC_1063 
+ TSMC_1064 TSMC_1065 TSMC_1066 TSMC_1067 TSMC_1068 TSMC_1069 
+ TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 TSMC_1074 TSMC_1075 
+ TSMC_1076 TSMC_1077 VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_537 
+ TSMC_538 TSMC_539 TSMC_540 TSMC_1057 TSMC_1058 
+ S1ALLSVTSW40W80_XDRV_LA512_884_SB 
XXDRV_LA512_SB_1 TSMC_1078 TSMC_1079 TSMC_1080 TSMC_1081 TSMC_1082 
+ TSMC_1083 TSMC_1084 TSMC_1085 TSMC_1067 TSMC_1086 TSMC_1087 
+ TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 TSMC_1092 TSMC_1093 
+ TSMC_1094 TSMC_1095 VDD VSS TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_541 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_1057 TSMC_1058 
+ S1ALLSVTSW40W80_XDRV_LA512_884_SB 
XXDRV_LA512_SB_2 TSMC_1059 TSMC_1060 TSMC_1061 TSMC_1062 TSMC_1096 
+ TSMC_1097 TSMC_1098 TSMC_1099 TSMC_1100 TSMC_1101 TSMC_1102 
+ TSMC_1103 TSMC_1104 TSMC_1105 TSMC_1106 TSMC_1107 TSMC_1108 
+ TSMC_1109 TSMC_1110 VDD VSS TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_1057 TSMC_1058 
+ S1ALLSVTSW40W80_XDRV_LA512_884_SB 
XXDRV_LA512_SB_3 TSMC_1078 TSMC_1079 TSMC_1080 TSMC_1081 TSMC_1111 
+ TSMC_1112 TSMC_1113 TSMC_1114 TSMC_1100 TSMC_1115 TSMC_1116 
+ TSMC_1117 TSMC_1118 TSMC_1119 TSMC_1120 TSMC_1121 TSMC_1122 
+ TSMC_1123 TSMC_1124 VDD VSS TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_549 
+ TSMC_550 TSMC_551 TSMC_552 TSMC_1057 TSMC_1058 
+ S1ALLSVTSW40W80_XDRV_LA512_884_SB 
XTRACKING_XB16X4 TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_569 TSMC_570 
+ TSMC_571 TSMC_572 TSMC_577 TSMC_578 TSMC_579 TSMC_580 TSMC_585 
+ TSMC_586 TSMC_587 TSMC_588 TSMC_593 TSMC_594 TSMC_595 TSMC_596 
+ TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_625 TSMC_626 
+ TSMC_627 TSMC_628 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_641 
+ TSMC_642 TSMC_643 TSMC_644 TSMC_649 TSMC_650 TSMC_651 TSMC_652 
+ TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_665 TSMC_666 TSMC_667 
+ TSMC_668 TSMC_673 TSMC_674 TSMC_675 TSMC_676 TSMC_681 TSMC_682 
+ TSMC_683 TSMC_684 TSMC_689 TSMC_690 TSMC_691 TSMC_692 TSMC_697 TSMC_698 
+ TSMC_699 TSMC_700 TSMC_705 TSMC_706 TSMC_707 TSMC_708 TSMC_713 
+ TSMC_714 TSMC_715 TSMC_716 TSMC_721 TSMC_722 TSMC_723 TSMC_724 
+ TSMC_729 TSMC_730 TSMC_731 TSMC_732 TSMC_737 TSMC_738 TSMC_739 
+ TSMC_740 TSMC_745 TSMC_746 TSMC_747 TSMC_748 TSMC_753 TSMC_754 
+ TSMC_755 TSMC_756 TSMC_761 TSMC_762 TSMC_763 TSMC_764 TSMC_769 
+ TSMC_770 TSMC_771 TSMC_772 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_785 TSMC_786 TSMC_787 TSMC_788 TSMC_793 TSMC_794 TSMC_795 
+ TSMC_796 TSMC_801 TSMC_802 TSMC_803 TSMC_804 TSMC_809 TSMC_810 
+ TSMC_811 TSMC_812 TSMC_817 TSMC_818 TSMC_819 TSMC_820 TSMC_825 TSMC_826 
+ TSMC_827 TSMC_828 TSMC_833 TSMC_834 TSMC_835 TSMC_836 TSMC_841 
+ TSMC_842 TSMC_843 TSMC_844 TSMC_849 TSMC_850 TSMC_851 TSMC_852 
+ TSMC_857 TSMC_858 TSMC_859 TSMC_860 TSMC_865 TSMC_866 TSMC_867 
+ TSMC_868 TSMC_873 TSMC_874 TSMC_875 TSMC_876 TSMC_881 TSMC_882 
+ TSMC_883 TSMC_884 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_897 
+ TSMC_898 TSMC_899 TSMC_900 TSMC_905 TSMC_906 TSMC_907 TSMC_908 
+ TSMC_913 TSMC_914 TSMC_915 TSMC_916 TSMC_921 TSMC_922 TSMC_923 
+ TSMC_924 TSMC_929 TSMC_930 TSMC_931 TSMC_932 TSMC_937 TSMC_938 
+ TSMC_939 TSMC_940 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_953 TSMC_954 
+ TSMC_955 TSMC_956 TSMC_961 TSMC_962 TSMC_963 TSMC_964 TSMC_969 
+ TSMC_970 TSMC_971 TSMC_972 TSMC_977 TSMC_978 TSMC_979 TSMC_980 
+ TSMC_985 TSMC_986 TSMC_987 TSMC_988 TSMC_993 TSMC_994 TSMC_995 
+ TSMC_996 TSMC_1001 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1009 
+ TSMC_1010 TSMC_1011 TSMC_1012 TSMC_1017 TSMC_1018 TSMC_1019 
+ TSMC_1020 TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1033 TSMC_1034 
+ TSMC_1035 TSMC_1036 TSMC_1041 TSMC_1042 TSMC_1043 TSMC_1044 
+ TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1125 VDD VDD VSS 
+ TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 
+ TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 
+ TSMC_551 TSMC_552 TSMC_1126 S1ALLSVTSW40W80_TRACKING_SB 
XMIOM4_L_0 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_1127 
+ BWEB[0] TSMC_1128 D[0] Q[0] TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 
+ TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 TSMC_1137 
+ S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_1 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_25 TSMC_26 TSMC_27 TSMC_28 
+ TSMC_1127 BWEB[1] TSMC_1128 D[1] Q[1] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_2 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_33 TSMC_34 TSMC_35 TSMC_36 
+ TSMC_1127 BWEB[2] TSMC_1128 D[2] Q[2] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_3 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_1127 BWEB[3] TSMC_1128 D[3] Q[3] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_4 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_1127 BWEB[4] TSMC_1128 D[4] Q[4] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_5 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_1127 BWEB[5] TSMC_1128 D[5] Q[5] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_6 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_1127 BWEB[6] TSMC_1128 D[6] Q[6] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_7 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_73 TSMC_74 TSMC_75 TSMC_76 
+ TSMC_1127 BWEB[7] TSMC_1128 D[7] Q[7] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_8 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_81 TSMC_82 TSMC_83 TSMC_84 
+ TSMC_1127 BWEB[8] TSMC_1128 D[8] Q[8] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_9 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_89 TSMC_90 TSMC_91 TSMC_92 
+ TSMC_1127 BWEB[9] TSMC_1128 D[9] Q[9] TSMC_1129 VDD VSS TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_10 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_97 TSMC_98 TSMC_99 
+ TSMC_100 TSMC_1127 BWEB[10] TSMC_1128 D[10] Q[10] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_11 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_105 TSMC_106 TSMC_107 
+ TSMC_108 TSMC_1127 BWEB[11] TSMC_1128 D[11] Q[11] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_12 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_113 TSMC_114 TSMC_115 
+ TSMC_116 TSMC_1127 BWEB[12] TSMC_1128 D[12] Q[12] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_13 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_1127 BWEB[13] TSMC_1128 D[13] Q[13] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_14 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_129 TSMC_130 TSMC_131 
+ TSMC_132 TSMC_1127 BWEB[14] TSMC_1128 D[14] Q[14] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_15 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_1127 BWEB[15] TSMC_1128 D[15] Q[15] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_16 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_145 TSMC_146 TSMC_147 
+ TSMC_148 TSMC_1127 BWEB[16] TSMC_1128 D[16] Q[16] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_17 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_153 TSMC_154 TSMC_155 
+ TSMC_156 TSMC_1127 BWEB[17] TSMC_1128 D[17] Q[17] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_18 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_161 TSMC_162 TSMC_163 
+ TSMC_164 TSMC_1127 BWEB[18] TSMC_1128 D[18] Q[18] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_19 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_169 TSMC_170 TSMC_171 
+ TSMC_172 TSMC_1127 BWEB[19] TSMC_1128 D[19] Q[19] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_20 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_1127 BWEB[20] TSMC_1128 D[20] Q[20] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_21 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_185 TSMC_186 TSMC_187 
+ TSMC_188 TSMC_1127 BWEB[21] TSMC_1128 D[21] Q[21] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_22 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_193 TSMC_194 TSMC_195 
+ TSMC_196 TSMC_1127 BWEB[22] TSMC_1128 D[22] Q[22] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_23 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_1127 BWEB[23] TSMC_1128 D[23] Q[23] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_24 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_1127 BWEB[24] TSMC_1128 D[24] Q[24] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_25 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_1127 BWEB[25] TSMC_1128 D[25] Q[25] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_26 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_225 TSMC_226 TSMC_227 
+ TSMC_228 TSMC_1127 BWEB[26] TSMC_1128 D[26] Q[26] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_27 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_1127 BWEB[27] TSMC_1128 D[27] Q[27] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_28 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_241 TSMC_242 TSMC_243 
+ TSMC_244 TSMC_1127 BWEB[28] TSMC_1128 D[28] Q[28] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_29 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_249 TSMC_250 TSMC_251 
+ TSMC_252 TSMC_1127 BWEB[29] TSMC_1128 D[29] Q[29] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_30 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_257 TSMC_258 TSMC_259 
+ TSMC_260 TSMC_1127 BWEB[30] TSMC_1128 D[30] Q[30] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_31 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_265 TSMC_266 TSMC_267 
+ TSMC_268 TSMC_1127 BWEB[31] TSMC_1128 D[31] Q[31] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_32 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_273 TSMC_274 TSMC_275 
+ TSMC_276 TSMC_1127 BWEB[32] TSMC_1128 D[32] Q[32] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_33 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_281 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_1127 BWEB[33] TSMC_1128 D[33] Q[33] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_34 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_289 TSMC_290 TSMC_291 
+ TSMC_292 TSMC_1127 BWEB[34] TSMC_1128 D[34] Q[34] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_35 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_297 TSMC_298 TSMC_299 
+ TSMC_300 TSMC_1127 BWEB[35] TSMC_1128 D[35] Q[35] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_36 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_305 TSMC_306 TSMC_307 
+ TSMC_308 TSMC_1127 BWEB[36] TSMC_1128 D[36] Q[36] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_37 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_313 TSMC_314 TSMC_315 
+ TSMC_316 TSMC_1127 BWEB[37] TSMC_1128 D[37] Q[37] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_38 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_321 TSMC_322 TSMC_323 
+ TSMC_324 TSMC_1127 BWEB[38] TSMC_1128 D[38] Q[38] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_39 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_329 TSMC_330 TSMC_331 
+ TSMC_332 TSMC_1127 BWEB[39] TSMC_1128 D[39] Q[39] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_40 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_1127 BWEB[40] TSMC_1128 D[40] Q[40] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_41 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_345 TSMC_346 TSMC_347 
+ TSMC_348 TSMC_1127 BWEB[41] TSMC_1128 D[41] Q[41] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_42 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_353 TSMC_354 TSMC_355 
+ TSMC_356 TSMC_1127 BWEB[42] TSMC_1128 D[42] Q[42] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_43 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_361 TSMC_362 TSMC_363 
+ TSMC_364 TSMC_1127 BWEB[43] TSMC_1128 D[43] Q[43] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_44 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_369 TSMC_370 TSMC_371 
+ TSMC_372 TSMC_1127 BWEB[44] TSMC_1128 D[44] Q[44] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_45 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_377 TSMC_378 TSMC_379 
+ TSMC_380 TSMC_1127 BWEB[45] TSMC_1128 D[45] Q[45] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_46 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_385 TSMC_386 TSMC_387 
+ TSMC_388 TSMC_1127 BWEB[46] TSMC_1128 D[46] Q[46] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_47 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_393 TSMC_394 TSMC_395 
+ TSMC_396 TSMC_1127 BWEB[47] TSMC_1128 D[47] Q[47] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_48 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_1127 BWEB[48] TSMC_1128 D[48] Q[48] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_49 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_1127 BWEB[49] TSMC_1128 D[49] Q[49] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_50 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_417 TSMC_418 TSMC_419 
+ TSMC_420 TSMC_1127 BWEB[50] TSMC_1128 D[50] Q[50] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_51 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_425 TSMC_426 TSMC_427 
+ TSMC_428 TSMC_1127 BWEB[51] TSMC_1128 D[51] Q[51] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_52 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_433 TSMC_434 TSMC_435 
+ TSMC_436 TSMC_1127 BWEB[52] TSMC_1128 D[52] Q[52] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_53 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_441 TSMC_442 TSMC_443 
+ TSMC_444 TSMC_1127 BWEB[53] TSMC_1128 D[53] Q[53] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_54 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_449 TSMC_450 TSMC_451 
+ TSMC_452 TSMC_1127 BWEB[54] TSMC_1128 D[54] Q[54] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_55 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_457 TSMC_458 TSMC_459 
+ TSMC_460 TSMC_1127 BWEB[55] TSMC_1128 D[55] Q[55] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_56 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_1127 BWEB[56] TSMC_1128 D[56] Q[56] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_57 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_1127 BWEB[57] TSMC_1128 D[57] Q[57] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_58 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_481 TSMC_482 TSMC_483 
+ TSMC_484 TSMC_1127 BWEB[58] TSMC_1128 D[58] Q[58] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_59 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_489 TSMC_490 TSMC_491 
+ TSMC_492 TSMC_1127 BWEB[59] TSMC_1128 D[59] Q[59] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_60 TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_497 TSMC_498 TSMC_499 
+ TSMC_500 TSMC_1127 BWEB[60] TSMC_1128 D[60] Q[60] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_61 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_505 TSMC_506 TSMC_507 
+ TSMC_508 TSMC_1127 BWEB[61] TSMC_1128 D[61] Q[61] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_62 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_513 TSMC_514 TSMC_515 
+ TSMC_516 TSMC_1127 BWEB[62] TSMC_1128 D[62] Q[62] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_L_63 TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_521 TSMC_522 TSMC_523 
+ TSMC_524 TSMC_1127 BWEB[63] TSMC_1128 D[63] Q[63] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_64 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_1138 BWEB[64] TSMC_1139 D[64] Q[64] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_65 TSMC_557 TSMC_558 TSMC_559 TSMC_560 TSMC_553 TSMC_554 TSMC_555 
+ TSMC_556 TSMC_1138 BWEB[65] TSMC_1139 D[65] Q[65] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_66 TSMC_565 TSMC_566 TSMC_567 TSMC_568 TSMC_561 TSMC_562 TSMC_563 
+ TSMC_564 TSMC_1138 BWEB[66] TSMC_1139 D[66] Q[66] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_67 TSMC_573 TSMC_574 TSMC_575 TSMC_576 TSMC_569 TSMC_570 TSMC_571 
+ TSMC_572 TSMC_1138 BWEB[67] TSMC_1139 D[67] Q[67] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_68 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_577 TSMC_578 TSMC_579 
+ TSMC_580 TSMC_1138 BWEB[68] TSMC_1139 D[68] Q[68] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_69 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_1138 BWEB[69] TSMC_1139 D[69] Q[69] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_70 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_593 TSMC_594 TSMC_595 
+ TSMC_596 TSMC_1138 BWEB[70] TSMC_1139 D[70] Q[70] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_71 TSMC_605 TSMC_606 TSMC_607 TSMC_608 TSMC_601 TSMC_602 TSMC_603 
+ TSMC_604 TSMC_1138 BWEB[71] TSMC_1139 D[71] Q[71] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_72 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_1138 BWEB[72] TSMC_1139 D[72] Q[72] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_73 TSMC_621 TSMC_622 TSMC_623 TSMC_624 TSMC_617 TSMC_618 TSMC_619 
+ TSMC_620 TSMC_1138 BWEB[73] TSMC_1139 D[73] Q[73] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_74 TSMC_629 TSMC_630 TSMC_631 TSMC_632 TSMC_625 TSMC_626 TSMC_627 
+ TSMC_628 TSMC_1138 BWEB[74] TSMC_1139 D[74] Q[74] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_75 TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_633 TSMC_634 TSMC_635 
+ TSMC_636 TSMC_1138 BWEB[75] TSMC_1139 D[75] Q[75] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_76 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_1138 BWEB[76] TSMC_1139 D[76] Q[76] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_77 TSMC_653 TSMC_654 TSMC_655 TSMC_656 TSMC_649 TSMC_650 TSMC_651 
+ TSMC_652 TSMC_1138 BWEB[77] TSMC_1139 D[77] Q[77] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_78 TSMC_661 TSMC_662 TSMC_663 TSMC_664 TSMC_657 TSMC_658 TSMC_659 
+ TSMC_660 TSMC_1138 BWEB[78] TSMC_1139 D[78] Q[78] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_79 TSMC_669 TSMC_670 TSMC_671 TSMC_672 TSMC_665 TSMC_666 TSMC_667 
+ TSMC_668 TSMC_1138 BWEB[79] TSMC_1139 D[79] Q[79] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_80 TSMC_677 TSMC_678 TSMC_679 TSMC_680 TSMC_673 TSMC_674 TSMC_675 
+ TSMC_676 TSMC_1138 BWEB[80] TSMC_1139 D[80] Q[80] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_81 TSMC_685 TSMC_686 TSMC_687 TSMC_688 TSMC_681 TSMC_682 TSMC_683 
+ TSMC_684 TSMC_1138 BWEB[81] TSMC_1139 D[81] Q[81] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_82 TSMC_693 TSMC_694 TSMC_695 TSMC_696 TSMC_689 TSMC_690 TSMC_691 
+ TSMC_692 TSMC_1138 BWEB[82] TSMC_1139 D[82] Q[82] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_83 TSMC_701 TSMC_702 TSMC_703 TSMC_704 TSMC_697 TSMC_698 TSMC_699 
+ TSMC_700 TSMC_1138 BWEB[83] TSMC_1139 D[83] Q[83] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_84 TSMC_709 TSMC_710 TSMC_711 TSMC_712 TSMC_705 TSMC_706 TSMC_707 
+ TSMC_708 TSMC_1138 BWEB[84] TSMC_1139 D[84] Q[84] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_85 TSMC_717 TSMC_718 TSMC_719 TSMC_720 TSMC_713 TSMC_714 TSMC_715 
+ TSMC_716 TSMC_1138 BWEB[85] TSMC_1139 D[85] Q[85] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_86 TSMC_725 TSMC_726 TSMC_727 TSMC_728 TSMC_721 TSMC_722 TSMC_723 
+ TSMC_724 TSMC_1138 BWEB[86] TSMC_1139 D[86] Q[86] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_87 TSMC_733 TSMC_734 TSMC_735 TSMC_736 TSMC_729 TSMC_730 TSMC_731 
+ TSMC_732 TSMC_1138 BWEB[87] TSMC_1139 D[87] Q[87] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_88 TSMC_741 TSMC_742 TSMC_743 TSMC_744 TSMC_737 TSMC_738 TSMC_739 
+ TSMC_740 TSMC_1138 BWEB[88] TSMC_1139 D[88] Q[88] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_89 TSMC_749 TSMC_750 TSMC_751 TSMC_752 TSMC_745 TSMC_746 TSMC_747 
+ TSMC_748 TSMC_1138 BWEB[89] TSMC_1139 D[89] Q[89] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_90 TSMC_757 TSMC_758 TSMC_759 TSMC_760 TSMC_753 TSMC_754 TSMC_755 
+ TSMC_756 TSMC_1138 BWEB[90] TSMC_1139 D[90] Q[90] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_91 TSMC_765 TSMC_766 TSMC_767 TSMC_768 TSMC_761 TSMC_762 TSMC_763 
+ TSMC_764 TSMC_1138 BWEB[91] TSMC_1139 D[91] Q[91] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_92 TSMC_773 TSMC_774 TSMC_775 TSMC_776 TSMC_769 TSMC_770 TSMC_771 
+ TSMC_772 TSMC_1138 BWEB[92] TSMC_1139 D[92] Q[92] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_93 TSMC_781 TSMC_782 TSMC_783 TSMC_784 TSMC_777 TSMC_778 TSMC_779 
+ TSMC_780 TSMC_1138 BWEB[93] TSMC_1139 D[93] Q[93] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_94 TSMC_789 TSMC_790 TSMC_791 TSMC_792 TSMC_785 TSMC_786 TSMC_787 
+ TSMC_788 TSMC_1138 BWEB[94] TSMC_1139 D[94] Q[94] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_95 TSMC_797 TSMC_798 TSMC_799 TSMC_800 TSMC_793 TSMC_794 TSMC_795 
+ TSMC_796 TSMC_1138 BWEB[95] TSMC_1139 D[95] Q[95] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_96 TSMC_805 TSMC_806 TSMC_807 TSMC_808 TSMC_801 TSMC_802 TSMC_803 
+ TSMC_804 TSMC_1138 BWEB[96] TSMC_1139 D[96] Q[96] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_97 TSMC_813 TSMC_814 TSMC_815 TSMC_816 TSMC_809 TSMC_810 TSMC_811 
+ TSMC_812 TSMC_1138 BWEB[97] TSMC_1139 D[97] Q[97] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_98 TSMC_821 TSMC_822 TSMC_823 TSMC_824 TSMC_817 TSMC_818 TSMC_819 
+ TSMC_820 TSMC_1138 BWEB[98] TSMC_1139 D[98] Q[98] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_99 TSMC_829 TSMC_830 TSMC_831 TSMC_832 TSMC_825 TSMC_826 TSMC_827 
+ TSMC_828 TSMC_1138 BWEB[99] TSMC_1139 D[99] Q[99] TSMC_1129 VDD VSS 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_100 TSMC_837 TSMC_838 TSMC_839 TSMC_840 TSMC_833 TSMC_834 TSMC_835 
+ TSMC_836 TSMC_1138 BWEB[100] TSMC_1139 D[100] Q[100] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_101 TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_841 TSMC_842 TSMC_843 
+ TSMC_844 TSMC_1138 BWEB[101] TSMC_1139 D[101] Q[101] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_102 TSMC_853 TSMC_854 TSMC_855 TSMC_856 TSMC_849 TSMC_850 TSMC_851 
+ TSMC_852 TSMC_1138 BWEB[102] TSMC_1139 D[102] Q[102] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_103 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_857 TSMC_858 TSMC_859 
+ TSMC_860 TSMC_1138 BWEB[103] TSMC_1139 D[103] Q[103] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_104 TSMC_869 TSMC_870 TSMC_871 TSMC_872 TSMC_865 TSMC_866 TSMC_867 
+ TSMC_868 TSMC_1138 BWEB[104] TSMC_1139 D[104] Q[104] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_105 TSMC_877 TSMC_878 TSMC_879 TSMC_880 TSMC_873 TSMC_874 TSMC_875 
+ TSMC_876 TSMC_1138 BWEB[105] TSMC_1139 D[105] Q[105] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_106 TSMC_885 TSMC_886 TSMC_887 TSMC_888 TSMC_881 TSMC_882 TSMC_883 
+ TSMC_884 TSMC_1138 BWEB[106] TSMC_1139 D[106] Q[106] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_107 TSMC_893 TSMC_894 TSMC_895 TSMC_896 TSMC_889 TSMC_890 TSMC_891 
+ TSMC_892 TSMC_1138 BWEB[107] TSMC_1139 D[107] Q[107] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_108 TSMC_901 TSMC_902 TSMC_903 TSMC_904 TSMC_897 TSMC_898 TSMC_899 
+ TSMC_900 TSMC_1138 BWEB[108] TSMC_1139 D[108] Q[108] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_109 TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_905 TSMC_906 TSMC_907 
+ TSMC_908 TSMC_1138 BWEB[109] TSMC_1139 D[109] Q[109] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_110 TSMC_917 TSMC_918 TSMC_919 TSMC_920 TSMC_913 TSMC_914 TSMC_915 
+ TSMC_916 TSMC_1138 BWEB[110] TSMC_1139 D[110] Q[110] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_111 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_921 TSMC_922 TSMC_923 
+ TSMC_924 TSMC_1138 BWEB[111] TSMC_1139 D[111] Q[111] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_112 TSMC_933 TSMC_934 TSMC_935 TSMC_936 TSMC_929 TSMC_930 TSMC_931 
+ TSMC_932 TSMC_1138 BWEB[112] TSMC_1139 D[112] Q[112] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_113 TSMC_941 TSMC_942 TSMC_943 TSMC_944 TSMC_937 TSMC_938 TSMC_939 
+ TSMC_940 TSMC_1138 BWEB[113] TSMC_1139 D[113] Q[113] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_114 TSMC_949 TSMC_950 TSMC_951 TSMC_952 TSMC_945 TSMC_946 TSMC_947 
+ TSMC_948 TSMC_1138 BWEB[114] TSMC_1139 D[114] Q[114] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_115 TSMC_957 TSMC_958 TSMC_959 TSMC_960 TSMC_953 TSMC_954 TSMC_955 
+ TSMC_956 TSMC_1138 BWEB[115] TSMC_1139 D[115] Q[115] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_116 TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_961 TSMC_962 TSMC_963 
+ TSMC_964 TSMC_1138 BWEB[116] TSMC_1139 D[116] Q[116] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_117 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_1138 BWEB[117] TSMC_1139 D[117] Q[117] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_118 TSMC_981 TSMC_982 TSMC_983 TSMC_984 TSMC_977 TSMC_978 TSMC_979 
+ TSMC_980 TSMC_1138 BWEB[118] TSMC_1139 D[118] Q[118] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_119 TSMC_989 TSMC_990 TSMC_991 TSMC_992 TSMC_985 TSMC_986 TSMC_987 
+ TSMC_988 TSMC_1138 BWEB[119] TSMC_1139 D[119] Q[119] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_120 TSMC_997 TSMC_998 TSMC_999 TSMC_1000 TSMC_993 TSMC_994 TSMC_995 
+ TSMC_996 TSMC_1138 BWEB[120] TSMC_1139 D[120] Q[120] TSMC_1129 VDD 
+ VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 
+ TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_121 TSMC_1005 TSMC_1006 TSMC_1007 TSMC_1008 TSMC_1001 TSMC_1002 
+ TSMC_1003 TSMC_1004 TSMC_1138 BWEB[121] TSMC_1139 D[121] Q[121] 
+ TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_122 TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1009 TSMC_1010 
+ TSMC_1011 TSMC_1012 TSMC_1138 BWEB[122] TSMC_1139 D[122] Q[122] 
+ TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_123 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1138 BWEB[123] TSMC_1139 D[123] Q[123] 
+ TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_124 TSMC_1029 TSMC_1030 TSMC_1031 TSMC_1032 TSMC_1025 TSMC_1026 
+ TSMC_1027 TSMC_1028 TSMC_1138 BWEB[124] TSMC_1139 D[124] Q[124] 
+ TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_125 TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1033 TSMC_1034 
+ TSMC_1035 TSMC_1036 TSMC_1138 BWEB[125] TSMC_1139 D[125] Q[125] 
+ TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_126 TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 TSMC_1041 TSMC_1042 
+ TSMC_1043 TSMC_1044 TSMC_1138 BWEB[126] TSMC_1139 D[126] Q[126] 
+ TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIOM4_R_127 TSMC_1053 TSMC_1054 TSMC_1055 TSMC_1056 TSMC_1049 TSMC_1050 
+ TSMC_1051 TSMC_1052 TSMC_1138 BWEB[127] TSMC_1139 D[127] Q[127] 
+ TSMC_1129 VDD VSS TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 S1ALLSVTSW40W80_MIO_SB 
XMIO_SB_EDGE_L VDD TSMC_1140 TSMC_1141 VSS 
+ S1ALLSVTSW40W80_MIO_SB_EDGE 
XMIO_SB_EDGE_R VDD TSMC_1140 TSMC_1141 VSS 
+ S1ALLSVTSW40W80_MIO_SB_EDGE 
XCNT_M4_SB TSMC_1127 TSMC_1138 TSMC_1126 CEB TSMC_1128 TSMC_1139 CLK TSMC_1059 
+ TSMC_1060 TSMC_1061 TSMC_1062 TSMC_1078 TSMC_1079 TSMC_1080 
+ TSMC_1081 TSMC_1067 TSMC_1100 TSMC_1142 TSMC_1143 TSMC_1144 
+ TSMC_1145 TSMC_1146 TSMC_1147 TSMC_1057 TSMC_1148 TSMC_1149 
+ TSMC_1150 TSMC_1151 TSMC_1152 TSMC_1153 TSMC_1154 TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 RTSEL[0] RTSEL[1] TSMC_1129 TSMC_1141 TSMC_1125 VDD VSS WEB 
+ WTSEL[0] WTSEL[1] TSMC_1141 A[2] A[3] A[4] A[5] TSMC_1141 TSMC_1141 
+ TSMC_1141 TSMC_1141 A[0] A[1] TSMC_1141 TSMC_1141 
+ S1ALLSVTSW40W80_CNT_M4_SB 
XD_WEB WEB TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_CEB CEB TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_CLK CLK TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_A0 A[0] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_A1 A[1] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_A2 A[2] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_A3 A[3] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_A4 A[4] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_A5 A[5] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_D0 D[0] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D1 D[1] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D2 D[2] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D3 D[3] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D4 D[4] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D5 D[5] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D6 D[6] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D7 D[7] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D8 D[8] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D9 D[9] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D10 D[10] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D11 D[11] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D12 D[12] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D13 D[13] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D14 D[14] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D15 D[15] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D16 D[16] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D17 D[17] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D18 D[18] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D19 D[19] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D20 D[20] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D21 D[21] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D22 D[22] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D23 D[23] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D24 D[24] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D25 D[25] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D26 D[26] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D27 D[27] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D28 D[28] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D29 D[29] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D30 D[30] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D31 D[31] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D32 D[32] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D33 D[33] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D34 D[34] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D35 D[35] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D36 D[36] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D37 D[37] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D38 D[38] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D39 D[39] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D40 D[40] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D41 D[41] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D42 D[42] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D43 D[43] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D44 D[44] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D45 D[45] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D46 D[46] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D47 D[47] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D48 D[48] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D49 D[49] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D50 D[50] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D51 D[51] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D52 D[52] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D53 D[53] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D54 D[54] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D55 D[55] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D56 D[56] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D57 D[57] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D58 D[58] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D59 D[59] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D60 D[60] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D61 D[61] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D62 D[62] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D63 D[63] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D64 D[64] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D65 D[65] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D66 D[66] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D67 D[67] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D68 D[68] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D69 D[69] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D70 D[70] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D71 D[71] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D72 D[72] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D73 D[73] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D74 D[74] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D75 D[75] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D76 D[76] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D77 D[77] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D78 D[78] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D79 D[79] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D80 D[80] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D81 D[81] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D82 D[82] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D83 D[83] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D84 D[84] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D85 D[85] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D86 D[86] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D87 D[87] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D88 D[88] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D89 D[89] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D90 D[90] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D91 D[91] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D92 D[92] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D93 D[93] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D94 D[94] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D95 D[95] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D96 D[96] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D97 D[97] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D98 D[98] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D99 D[99] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D100 D[100] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D101 D[101] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D102 D[102] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D103 D[103] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D104 D[104] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D105 D[105] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D106 D[106] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D107 D[107] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D108 D[108] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D109 D[109] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D110 D[110] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D111 D[111] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D112 D[112] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D113 D[113] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D114 D[114] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D115 D[115] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D116 D[116] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D117 D[117] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D118 D[118] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D119 D[119] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D120 D[120] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D121 D[121] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D122 D[122] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D123 D[123] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D124 D[124] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D125 D[125] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D126 D[126] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_D127 D[127] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB0 BWEB[0] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB1 BWEB[1] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB2 BWEB[2] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB3 BWEB[3] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB4 BWEB[4] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB5 BWEB[5] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB6 BWEB[6] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB7 BWEB[7] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB8 BWEB[8] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB9 BWEB[9] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB10 BWEB[10] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB11 BWEB[11] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB12 BWEB[12] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB13 BWEB[13] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB14 BWEB[14] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB15 BWEB[15] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB16 BWEB[16] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB17 BWEB[17] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB18 BWEB[18] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB19 BWEB[19] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB20 BWEB[20] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB21 BWEB[21] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB22 BWEB[22] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB23 BWEB[23] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB24 BWEB[24] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB25 BWEB[25] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB26 BWEB[26] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB27 BWEB[27] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB28 BWEB[28] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB29 BWEB[29] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB30 BWEB[30] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB31 BWEB[31] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB32 BWEB[32] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB33 BWEB[33] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB34 BWEB[34] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB35 BWEB[35] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB36 BWEB[36] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB37 BWEB[37] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB38 BWEB[38] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB39 BWEB[39] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB40 BWEB[40] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB41 BWEB[41] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB42 BWEB[42] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB43 BWEB[43] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB44 BWEB[44] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB45 BWEB[45] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB46 BWEB[46] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB47 BWEB[47] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB48 BWEB[48] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB49 BWEB[49] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB50 BWEB[50] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB51 BWEB[51] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB52 BWEB[52] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB53 BWEB[53] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB54 BWEB[54] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB55 BWEB[55] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB56 BWEB[56] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB57 BWEB[57] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB58 BWEB[58] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB59 BWEB[59] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB60 BWEB[60] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB61 BWEB[61] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB62 BWEB[62] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB63 BWEB[63] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB64 BWEB[64] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB65 BWEB[65] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB66 BWEB[66] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB67 BWEB[67] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB68 BWEB[68] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB69 BWEB[69] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB70 BWEB[70] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB71 BWEB[71] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB72 BWEB[72] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB73 BWEB[73] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB74 BWEB[74] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB75 BWEB[75] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB76 BWEB[76] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB77 BWEB[77] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB78 BWEB[78] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB79 BWEB[79] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB80 BWEB[80] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB81 BWEB[81] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB82 BWEB[82] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB83 BWEB[83] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB84 BWEB[84] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB85 BWEB[85] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB86 BWEB[86] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB87 BWEB[87] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB88 BWEB[88] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB89 BWEB[89] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB90 BWEB[90] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB91 BWEB[91] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB92 BWEB[92] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB93 BWEB[93] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB94 BWEB[94] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB95 BWEB[95] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB96 BWEB[96] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB97 BWEB[97] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB98 BWEB[98] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB99 BWEB[99] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB100 BWEB[100] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB101 BWEB[101] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB102 BWEB[102] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB103 BWEB[103] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB104 BWEB[104] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB105 BWEB[105] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB106 BWEB[106] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB107 BWEB[107] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB108 BWEB[108] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB109 BWEB[109] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB110 BWEB[110] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB111 BWEB[111] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB112 BWEB[112] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB113 BWEB[113] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB114 BWEB[114] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB115 BWEB[115] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB116 BWEB[116] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB117 BWEB[117] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB118 BWEB[118] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB119 BWEB[119] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB120 BWEB[120] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB121 BWEB[121] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB122 BWEB[122] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB123 BWEB[123] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB124 BWEB[124] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB125 BWEB[125] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB126 BWEB[126] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_BWEB127 BWEB[127] VSS S1ALLSVTSW40W80_DIO_TALL 
XD_WTESL_1 WTSEL[1] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_WTESL_0 WTSEL[0] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_RTESL_1 RTSEL[1] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
XD_RTESL_0 RTSEL[0] TSMC_1141 VSS S1ALLSVTSW40W80_DIODE 
.ENDS


