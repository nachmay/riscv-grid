# Created by MC2 : Version 2013.12.00.f on 2025/06/18, 12:43:53

 
###############################################################################
#                                                    
#        Technology     : TSMC 16nm CMOS Logic FinFet (FFC) HKMG
#        Memory Type    : TSMC 16nm FFC Two Port Register File with d130 bit cell
#        Library Name   : ts6n16ffcllsvta32x32m4fw (user specify : ts6n16ffcllsvta32x32m4fw)
#        Library Version: 170a
#        Generated Time : 2025/06/18, 12:42:56
###############################################################################
# STATEMENT OF USE                                                             
#                                                                              
#  This information contains confidential and proprietary information of TSMC. 
# No part of this information may be reproduced, transmitted, transcribed,     
# stored in a retrieval system, or translated into any human or computer       
# language, in any form or by any means, electronic, mechanical, magnetic,     
# optical, chemical, manual, or otherwise, without the prior written permission
# of TSMC. This information was prepared for informational purpose and is for  
# use by TSMC's customers only. TSMC reserves the right to make changes in the 
# inforrmation at any time and without notice.                                 
###############################################################################
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
#                                                                              

MACRO TS6N16FFCLLSVTA32X32M4FW
	CLASS BLOCK ;
	FOREIGN TS6N16FFCLLSVTA32X32M4FW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 15.517 BY 112.800 ;
	SYMMETRY X Y ;
	PIN AA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 52.142 15.517 52.222 ;
			LAYER M2 ;
			RECT 15.269 52.142 15.517 52.222 ;
			LAYER M3 ;
			RECT 15.269 52.142 15.517 52.222 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[0]

	PIN AA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 52.370 15.517 52.450 ;
			LAYER M2 ;
			RECT 15.269 52.370 15.517 52.450 ;
			LAYER M3 ;
			RECT 15.269 52.370 15.517 52.450 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[1]

	PIN AA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 55.334 15.517 55.414 ;
			LAYER M2 ;
			RECT 15.269 55.334 15.517 55.414 ;
			LAYER M3 ;
			RECT 15.269 55.334 15.517 55.414 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[2]

	PIN AA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 53.738 15.517 53.818 ;
			LAYER M2 ;
			RECT 15.269 53.738 15.517 53.818 ;
			LAYER M3 ;
			RECT 15.269 53.738 15.517 53.818 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[3]

	PIN AA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 55.106 15.517 55.186 ;
			LAYER M2 ;
			RECT 15.269 55.106 15.517 55.186 ;
			LAYER M3 ;
			RECT 15.269 55.106 15.517 55.186 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[4]

	PIN AB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 60.578 15.517 60.658 ;
			LAYER M2 ;
			RECT 15.269 60.578 15.517 60.658 ;
			LAYER M3 ;
			RECT 15.269 60.578 15.517 60.658 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[0]

	PIN AB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 60.350 15.517 60.430 ;
			LAYER M2 ;
			RECT 15.269 60.350 15.517 60.430 ;
			LAYER M3 ;
			RECT 15.269 60.350 15.517 60.430 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[1]

	PIN AB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 57.386 15.517 57.466 ;
			LAYER M2 ;
			RECT 15.269 57.386 15.517 57.466 ;
			LAYER M3 ;
			RECT 15.269 57.386 15.517 57.466 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[2]

	PIN AB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 58.982 15.517 59.062 ;
			LAYER M2 ;
			RECT 15.269 58.982 15.517 59.062 ;
			LAYER M3 ;
			RECT 15.269 58.982 15.517 59.062 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[3]

	PIN AB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 57.614 15.517 57.694 ;
			LAYER M2 ;
			RECT 15.269 57.614 15.517 57.694 ;
			LAYER M3 ;
			RECT 15.269 57.614 15.517 57.694 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[4]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 1.799 15.517 1.879 ;
			LAYER M2 ;
			RECT 15.269 1.799 15.517 1.879 ;
			LAYER M3 ;
			RECT 15.269 1.799 15.517 1.879 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 4.679 15.517 4.759 ;
			LAYER M2 ;
			RECT 15.269 4.679 15.517 4.759 ;
			LAYER M3 ;
			RECT 15.269 4.679 15.517 4.759 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 7.559 15.517 7.639 ;
			LAYER M2 ;
			RECT 15.269 7.559 15.517 7.639 ;
			LAYER M3 ;
			RECT 15.269 7.559 15.517 7.639 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 10.439 15.517 10.519 ;
			LAYER M2 ;
			RECT 15.269 10.439 15.517 10.519 ;
			LAYER M3 ;
			RECT 15.269 10.439 15.517 10.519 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 13.319 15.517 13.399 ;
			LAYER M2 ;
			RECT 15.269 13.319 15.517 13.399 ;
			LAYER M3 ;
			RECT 15.269 13.319 15.517 13.399 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 16.199 15.517 16.279 ;
			LAYER M2 ;
			RECT 15.269 16.199 15.517 16.279 ;
			LAYER M3 ;
			RECT 15.269 16.199 15.517 16.279 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 19.079 15.517 19.159 ;
			LAYER M2 ;
			RECT 15.269 19.079 15.517 19.159 ;
			LAYER M3 ;
			RECT 15.269 19.079 15.517 19.159 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 21.959 15.517 22.039 ;
			LAYER M2 ;
			RECT 15.269 21.959 15.517 22.039 ;
			LAYER M3 ;
			RECT 15.269 21.959 15.517 22.039 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 24.839 15.517 24.919 ;
			LAYER M2 ;
			RECT 15.269 24.839 15.517 24.919 ;
			LAYER M3 ;
			RECT 15.269 24.839 15.517 24.919 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 27.719 15.517 27.799 ;
			LAYER M2 ;
			RECT 15.269 27.719 15.517 27.799 ;
			LAYER M3 ;
			RECT 15.269 27.719 15.517 27.799 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 30.599 15.517 30.679 ;
			LAYER M2 ;
			RECT 15.269 30.599 15.517 30.679 ;
			LAYER M3 ;
			RECT 15.269 30.599 15.517 30.679 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 33.479 15.517 33.559 ;
			LAYER M2 ;
			RECT 15.269 33.479 15.517 33.559 ;
			LAYER M3 ;
			RECT 15.269 33.479 15.517 33.559 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 36.359 15.517 36.439 ;
			LAYER M2 ;
			RECT 15.269 36.359 15.517 36.439 ;
			LAYER M3 ;
			RECT 15.269 36.359 15.517 36.439 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 39.239 15.517 39.319 ;
			LAYER M2 ;
			RECT 15.269 39.239 15.517 39.319 ;
			LAYER M3 ;
			RECT 15.269 39.239 15.517 39.319 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 42.119 15.517 42.199 ;
			LAYER M2 ;
			RECT 15.269 42.119 15.517 42.199 ;
			LAYER M3 ;
			RECT 15.269 42.119 15.517 42.199 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 44.999 15.517 45.079 ;
			LAYER M2 ;
			RECT 15.269 44.999 15.517 45.079 ;
			LAYER M3 ;
			RECT 15.269 44.999 15.517 45.079 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 67.721 15.517 67.801 ;
			LAYER M2 ;
			RECT 15.269 67.721 15.517 67.801 ;
			LAYER M3 ;
			RECT 15.269 67.721 15.517 67.801 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 70.601 15.517 70.681 ;
			LAYER M2 ;
			RECT 15.269 70.601 15.517 70.681 ;
			LAYER M3 ;
			RECT 15.269 70.601 15.517 70.681 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 73.481 15.517 73.561 ;
			LAYER M2 ;
			RECT 15.269 73.481 15.517 73.561 ;
			LAYER M3 ;
			RECT 15.269 73.481 15.517 73.561 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 76.361 15.517 76.441 ;
			LAYER M2 ;
			RECT 15.269 76.361 15.517 76.441 ;
			LAYER M3 ;
			RECT 15.269 76.361 15.517 76.441 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 79.241 15.517 79.321 ;
			LAYER M2 ;
			RECT 15.269 79.241 15.517 79.321 ;
			LAYER M3 ;
			RECT 15.269 79.241 15.517 79.321 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 82.121 15.517 82.201 ;
			LAYER M2 ;
			RECT 15.269 82.121 15.517 82.201 ;
			LAYER M3 ;
			RECT 15.269 82.121 15.517 82.201 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 85.001 15.517 85.081 ;
			LAYER M2 ;
			RECT 15.269 85.001 15.517 85.081 ;
			LAYER M3 ;
			RECT 15.269 85.001 15.517 85.081 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 87.881 15.517 87.961 ;
			LAYER M2 ;
			RECT 15.269 87.881 15.517 87.961 ;
			LAYER M3 ;
			RECT 15.269 87.881 15.517 87.961 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 90.761 15.517 90.841 ;
			LAYER M2 ;
			RECT 15.269 90.761 15.517 90.841 ;
			LAYER M3 ;
			RECT 15.269 90.761 15.517 90.841 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 93.641 15.517 93.721 ;
			LAYER M2 ;
			RECT 15.269 93.641 15.517 93.721 ;
			LAYER M3 ;
			RECT 15.269 93.641 15.517 93.721 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 96.521 15.517 96.601 ;
			LAYER M2 ;
			RECT 15.269 96.521 15.517 96.601 ;
			LAYER M3 ;
			RECT 15.269 96.521 15.517 96.601 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 99.401 15.517 99.481 ;
			LAYER M2 ;
			RECT 15.269 99.401 15.517 99.481 ;
			LAYER M3 ;
			RECT 15.269 99.401 15.517 99.481 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 102.281 15.517 102.361 ;
			LAYER M2 ;
			RECT 15.269 102.281 15.517 102.361 ;
			LAYER M3 ;
			RECT 15.269 102.281 15.517 102.361 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 105.161 15.517 105.241 ;
			LAYER M2 ;
			RECT 15.269 105.161 15.517 105.241 ;
			LAYER M3 ;
			RECT 15.269 105.161 15.517 105.241 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 108.041 15.517 108.121 ;
			LAYER M2 ;
			RECT 15.269 108.041 15.517 108.121 ;
			LAYER M3 ;
			RECT 15.269 108.041 15.517 108.121 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 110.921 15.517 111.001 ;
			LAYER M2 ;
			RECT 15.269 110.921 15.517 111.001 ;
			LAYER M3 ;
			RECT 15.269 110.921 15.517 111.001 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[31]

	PIN CLKR
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 63.314 15.517 63.394 ;
			LAYER M2 ;
			RECT 15.269 63.314 15.517 63.394 ;
			LAYER M3 ;
			RECT 15.269 63.314 15.517 63.394 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2280 LAYER M2 ;
		ANTENNAMAXAREACAR 40.1766 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0128 LAYER M3 ;
		ANTENNAMAXAREACAR 179.9160 LAYER M3 ;
	END CLKR

	PIN CLKW
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 48.722 15.517 48.802 ;
			LAYER M2 ;
			RECT 15.269 48.722 15.517 48.802 ;
			LAYER M3 ;
			RECT 15.269 48.722 15.517 48.802 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.4639 LAYER M2 ;
		ANTENNAMAXAREACAR 44.8112 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0082 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0159 LAYER M3 ;
		ANTENNAMAXAREACAR 150.9920 LAYER M3 ;
	END CLKW

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 2.951 15.517 3.031 ;
			LAYER M2 ;
			RECT 15.269 2.951 15.517 3.031 ;
			LAYER M3 ;
			RECT 15.269 2.951 15.517 3.031 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 5.831 15.517 5.911 ;
			LAYER M2 ;
			RECT 15.269 5.831 15.517 5.911 ;
			LAYER M3 ;
			RECT 15.269 5.831 15.517 5.911 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 8.711 15.517 8.791 ;
			LAYER M2 ;
			RECT 15.269 8.711 15.517 8.791 ;
			LAYER M3 ;
			RECT 15.269 8.711 15.517 8.791 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 11.591 15.517 11.671 ;
			LAYER M2 ;
			RECT 15.269 11.591 15.517 11.671 ;
			LAYER M3 ;
			RECT 15.269 11.591 15.517 11.671 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 14.471 15.517 14.551 ;
			LAYER M2 ;
			RECT 15.269 14.471 15.517 14.551 ;
			LAYER M3 ;
			RECT 15.269 14.471 15.517 14.551 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 17.351 15.517 17.431 ;
			LAYER M2 ;
			RECT 15.269 17.351 15.517 17.431 ;
			LAYER M3 ;
			RECT 15.269 17.351 15.517 17.431 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 20.231 15.517 20.311 ;
			LAYER M2 ;
			RECT 15.269 20.231 15.517 20.311 ;
			LAYER M3 ;
			RECT 15.269 20.231 15.517 20.311 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 23.111 15.517 23.191 ;
			LAYER M2 ;
			RECT 15.269 23.111 15.517 23.191 ;
			LAYER M3 ;
			RECT 15.269 23.111 15.517 23.191 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 25.991 15.517 26.071 ;
			LAYER M2 ;
			RECT 15.269 25.991 15.517 26.071 ;
			LAYER M3 ;
			RECT 15.269 25.991 15.517 26.071 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 28.871 15.517 28.951 ;
			LAYER M2 ;
			RECT 15.269 28.871 15.517 28.951 ;
			LAYER M3 ;
			RECT 15.269 28.871 15.517 28.951 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 31.751 15.517 31.831 ;
			LAYER M2 ;
			RECT 15.269 31.751 15.517 31.831 ;
			LAYER M3 ;
			RECT 15.269 31.751 15.517 31.831 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 34.631 15.517 34.711 ;
			LAYER M2 ;
			RECT 15.269 34.631 15.517 34.711 ;
			LAYER M3 ;
			RECT 15.269 34.631 15.517 34.711 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 37.511 15.517 37.591 ;
			LAYER M2 ;
			RECT 15.269 37.511 15.517 37.591 ;
			LAYER M3 ;
			RECT 15.269 37.511 15.517 37.591 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 40.391 15.517 40.471 ;
			LAYER M2 ;
			RECT 15.269 40.391 15.517 40.471 ;
			LAYER M3 ;
			RECT 15.269 40.391 15.517 40.471 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 43.271 15.517 43.351 ;
			LAYER M2 ;
			RECT 15.269 43.271 15.517 43.351 ;
			LAYER M3 ;
			RECT 15.269 43.271 15.517 43.351 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 46.151 15.517 46.231 ;
			LAYER M2 ;
			RECT 15.269 46.151 15.517 46.231 ;
			LAYER M3 ;
			RECT 15.269 46.151 15.517 46.231 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 66.569 15.517 66.649 ;
			LAYER M2 ;
			RECT 15.269 66.569 15.517 66.649 ;
			LAYER M3 ;
			RECT 15.269 66.569 15.517 66.649 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 69.449 15.517 69.529 ;
			LAYER M2 ;
			RECT 15.269 69.449 15.517 69.529 ;
			LAYER M3 ;
			RECT 15.269 69.449 15.517 69.529 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 72.329 15.517 72.409 ;
			LAYER M2 ;
			RECT 15.269 72.329 15.517 72.409 ;
			LAYER M3 ;
			RECT 15.269 72.329 15.517 72.409 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 75.209 15.517 75.289 ;
			LAYER M2 ;
			RECT 15.269 75.209 15.517 75.289 ;
			LAYER M3 ;
			RECT 15.269 75.209 15.517 75.289 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 78.089 15.517 78.169 ;
			LAYER M2 ;
			RECT 15.269 78.089 15.517 78.169 ;
			LAYER M3 ;
			RECT 15.269 78.089 15.517 78.169 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 80.969 15.517 81.049 ;
			LAYER M2 ;
			RECT 15.269 80.969 15.517 81.049 ;
			LAYER M3 ;
			RECT 15.269 80.969 15.517 81.049 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 83.849 15.517 83.929 ;
			LAYER M2 ;
			RECT 15.269 83.849 15.517 83.929 ;
			LAYER M3 ;
			RECT 15.269 83.849 15.517 83.929 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 86.729 15.517 86.809 ;
			LAYER M2 ;
			RECT 15.269 86.729 15.517 86.809 ;
			LAYER M3 ;
			RECT 15.269 86.729 15.517 86.809 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 89.609 15.517 89.689 ;
			LAYER M2 ;
			RECT 15.269 89.609 15.517 89.689 ;
			LAYER M3 ;
			RECT 15.269 89.609 15.517 89.689 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 92.489 15.517 92.569 ;
			LAYER M2 ;
			RECT 15.269 92.489 15.517 92.569 ;
			LAYER M3 ;
			RECT 15.269 92.489 15.517 92.569 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 95.369 15.517 95.449 ;
			LAYER M2 ;
			RECT 15.269 95.369 15.517 95.449 ;
			LAYER M3 ;
			RECT 15.269 95.369 15.517 95.449 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 98.249 15.517 98.329 ;
			LAYER M2 ;
			RECT 15.269 98.249 15.517 98.329 ;
			LAYER M3 ;
			RECT 15.269 98.249 15.517 98.329 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 101.129 15.517 101.209 ;
			LAYER M2 ;
			RECT 15.269 101.129 15.517 101.209 ;
			LAYER M3 ;
			RECT 15.269 101.129 15.517 101.209 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 104.009 15.517 104.089 ;
			LAYER M2 ;
			RECT 15.269 104.009 15.517 104.089 ;
			LAYER M3 ;
			RECT 15.269 104.009 15.517 104.089 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 106.889 15.517 106.969 ;
			LAYER M2 ;
			RECT 15.269 106.889 15.517 106.969 ;
			LAYER M3 ;
			RECT 15.269 106.889 15.517 106.969 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 109.769 15.517 109.849 ;
			LAYER M2 ;
			RECT 15.269 109.769 15.517 109.849 ;
			LAYER M3 ;
			RECT 15.269 109.769 15.517 109.849 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[31]

	PIN KP[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 50.090 15.517 50.170 ;
			LAYER M2 ;
			RECT 15.269 50.090 15.517 50.170 ;
			LAYER M3 ;
			RECT 15.269 50.090 15.517 50.170 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[0]

	PIN KP[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 50.318 15.517 50.398 ;
			LAYER M2 ;
			RECT 15.269 50.318 15.517 50.398 ;
			LAYER M3 ;
			RECT 15.269 50.318 15.517 50.398 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[1]

	PIN KP[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 50.546 15.517 50.626 ;
			LAYER M2 ;
			RECT 15.269 50.546 15.517 50.626 ;
			LAYER M3 ;
			RECT 15.269 50.546 15.517 50.626 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[2]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 2.375 15.517 2.455 ;
			LAYER M2 ;
			RECT 15.269 2.375 15.517 2.455 ;
			LAYER M3 ;
			RECT 15.269 2.375 15.517 2.455 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 5.255 15.517 5.335 ;
			LAYER M2 ;
			RECT 15.269 5.255 15.517 5.335 ;
			LAYER M3 ;
			RECT 15.269 5.255 15.517 5.335 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 8.135 15.517 8.215 ;
			LAYER M2 ;
			RECT 15.269 8.135 15.517 8.215 ;
			LAYER M3 ;
			RECT 15.269 8.135 15.517 8.215 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 11.015 15.517 11.095 ;
			LAYER M2 ;
			RECT 15.269 11.015 15.517 11.095 ;
			LAYER M3 ;
			RECT 15.269 11.015 15.517 11.095 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 13.895 15.517 13.975 ;
			LAYER M2 ;
			RECT 15.269 13.895 15.517 13.975 ;
			LAYER M3 ;
			RECT 15.269 13.895 15.517 13.975 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 16.775 15.517 16.855 ;
			LAYER M2 ;
			RECT 15.269 16.775 15.517 16.855 ;
			LAYER M3 ;
			RECT 15.269 16.775 15.517 16.855 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 19.655 15.517 19.735 ;
			LAYER M2 ;
			RECT 15.269 19.655 15.517 19.735 ;
			LAYER M3 ;
			RECT 15.269 19.655 15.517 19.735 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 22.535 15.517 22.615 ;
			LAYER M2 ;
			RECT 15.269 22.535 15.517 22.615 ;
			LAYER M3 ;
			RECT 15.269 22.535 15.517 22.615 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 25.415 15.517 25.495 ;
			LAYER M2 ;
			RECT 15.269 25.415 15.517 25.495 ;
			LAYER M3 ;
			RECT 15.269 25.415 15.517 25.495 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 28.295 15.517 28.375 ;
			LAYER M2 ;
			RECT 15.269 28.295 15.517 28.375 ;
			LAYER M3 ;
			RECT 15.269 28.295 15.517 28.375 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 31.175 15.517 31.255 ;
			LAYER M2 ;
			RECT 15.269 31.175 15.517 31.255 ;
			LAYER M3 ;
			RECT 15.269 31.175 15.517 31.255 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 34.055 15.517 34.135 ;
			LAYER M2 ;
			RECT 15.269 34.055 15.517 34.135 ;
			LAYER M3 ;
			RECT 15.269 34.055 15.517 34.135 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 36.935 15.517 37.015 ;
			LAYER M2 ;
			RECT 15.269 36.935 15.517 37.015 ;
			LAYER M3 ;
			RECT 15.269 36.935 15.517 37.015 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 39.815 15.517 39.895 ;
			LAYER M2 ;
			RECT 15.269 39.815 15.517 39.895 ;
			LAYER M3 ;
			RECT 15.269 39.815 15.517 39.895 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 42.695 15.517 42.775 ;
			LAYER M2 ;
			RECT 15.269 42.695 15.517 42.775 ;
			LAYER M3 ;
			RECT 15.269 42.695 15.517 42.775 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 45.575 15.517 45.655 ;
			LAYER M2 ;
			RECT 15.269 45.575 15.517 45.655 ;
			LAYER M3 ;
			RECT 15.269 45.575 15.517 45.655 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 67.145 15.517 67.225 ;
			LAYER M2 ;
			RECT 15.269 67.145 15.517 67.225 ;
			LAYER M3 ;
			RECT 15.269 67.145 15.517 67.225 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 70.025 15.517 70.105 ;
			LAYER M2 ;
			RECT 15.269 70.025 15.517 70.105 ;
			LAYER M3 ;
			RECT 15.269 70.025 15.517 70.105 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 72.905 15.517 72.985 ;
			LAYER M2 ;
			RECT 15.269 72.905 15.517 72.985 ;
			LAYER M3 ;
			RECT 15.269 72.905 15.517 72.985 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 75.785 15.517 75.865 ;
			LAYER M2 ;
			RECT 15.269 75.785 15.517 75.865 ;
			LAYER M3 ;
			RECT 15.269 75.785 15.517 75.865 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 78.665 15.517 78.745 ;
			LAYER M2 ;
			RECT 15.269 78.665 15.517 78.745 ;
			LAYER M3 ;
			RECT 15.269 78.665 15.517 78.745 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 81.545 15.517 81.625 ;
			LAYER M2 ;
			RECT 15.269 81.545 15.517 81.625 ;
			LAYER M3 ;
			RECT 15.269 81.545 15.517 81.625 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 84.425 15.517 84.505 ;
			LAYER M2 ;
			RECT 15.269 84.425 15.517 84.505 ;
			LAYER M3 ;
			RECT 15.269 84.425 15.517 84.505 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 87.305 15.517 87.385 ;
			LAYER M2 ;
			RECT 15.269 87.305 15.517 87.385 ;
			LAYER M3 ;
			RECT 15.269 87.305 15.517 87.385 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 90.185 15.517 90.265 ;
			LAYER M2 ;
			RECT 15.269 90.185 15.517 90.265 ;
			LAYER M3 ;
			RECT 15.269 90.185 15.517 90.265 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 93.065 15.517 93.145 ;
			LAYER M2 ;
			RECT 15.269 93.065 15.517 93.145 ;
			LAYER M3 ;
			RECT 15.269 93.065 15.517 93.145 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 95.945 15.517 96.025 ;
			LAYER M2 ;
			RECT 15.269 95.945 15.517 96.025 ;
			LAYER M3 ;
			RECT 15.269 95.945 15.517 96.025 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 98.825 15.517 98.905 ;
			LAYER M2 ;
			RECT 15.269 98.825 15.517 98.905 ;
			LAYER M3 ;
			RECT 15.269 98.825 15.517 98.905 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 101.705 15.517 101.785 ;
			LAYER M2 ;
			RECT 15.269 101.705 15.517 101.785 ;
			LAYER M3 ;
			RECT 15.269 101.705 15.517 101.785 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 104.585 15.517 104.665 ;
			LAYER M2 ;
			RECT 15.269 104.585 15.517 104.665 ;
			LAYER M3 ;
			RECT 15.269 104.585 15.517 104.665 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 107.465 15.517 107.545 ;
			LAYER M2 ;
			RECT 15.269 107.465 15.517 107.545 ;
			LAYER M3 ;
			RECT 15.269 107.465 15.517 107.545 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 110.345 15.517 110.425 ;
			LAYER M2 ;
			RECT 15.269 110.345 15.517 110.425 ;
			LAYER M3 ;
			RECT 15.269 110.345 15.517 110.425 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[31]

	PIN RCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 65.138 15.517 65.218 ;
			LAYER M2 ;
			RECT 15.269 65.138 15.517 65.218 ;
			LAYER M3 ;
			RECT 15.269 65.138 15.517 65.218 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[0]

	PIN RCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 64.910 15.517 64.990 ;
			LAYER M2 ;
			RECT 15.269 64.910 15.517 64.990 ;
			LAYER M3 ;
			RECT 15.269 64.910 15.517 64.990 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[1]

	PIN REB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 61.490 15.517 61.570 ;
			LAYER M2 ;
			RECT 15.269 61.490 15.517 61.570 ;
			LAYER M3 ;
			RECT 15.269 61.490 15.517 61.570 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0860 LAYER M1 ;
		ANTENNAMAXAREACAR 12.8828 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0840 LAYER M2 ;
		ANTENNAMAXAREACAR 20.5069 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4602 LAYER M3 ;
		ANTENNAMAXAREACAR 218.8550 LAYER M3 ;
	END REB

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.624 15.397 1.784 ;
			LAYER M4 ;
			RECT 0.120 3.064 15.397 3.224 ;
			LAYER M4 ;
			RECT 0.120 4.504 15.397 4.664 ;
			LAYER M4 ;
			RECT 0.120 5.944 15.397 6.104 ;
			LAYER M4 ;
			RECT 0.120 7.384 15.397 7.544 ;
			LAYER M4 ;
			RECT 0.120 8.824 15.397 8.984 ;
			LAYER M4 ;
			RECT 0.120 10.264 15.397 10.424 ;
			LAYER M4 ;
			RECT 0.120 11.704 15.397 11.864 ;
			LAYER M4 ;
			RECT 0.120 13.144 15.397 13.304 ;
			LAYER M4 ;
			RECT 0.120 14.584 15.397 14.744 ;
			LAYER M4 ;
			RECT 0.120 16.024 15.397 16.184 ;
			LAYER M4 ;
			RECT 0.120 17.464 15.397 17.624 ;
			LAYER M4 ;
			RECT 0.120 18.904 15.397 19.064 ;
			LAYER M4 ;
			RECT 0.120 20.344 15.397 20.504 ;
			LAYER M4 ;
			RECT 0.120 21.784 15.397 21.944 ;
			LAYER M4 ;
			RECT 0.120 23.224 15.397 23.384 ;
			LAYER M4 ;
			RECT 0.120 24.664 15.397 24.824 ;
			LAYER M4 ;
			RECT 0.120 26.104 15.397 26.264 ;
			LAYER M4 ;
			RECT 0.120 27.544 15.397 27.704 ;
			LAYER M4 ;
			RECT 0.120 28.984 15.397 29.144 ;
			LAYER M4 ;
			RECT 0.120 30.424 15.397 30.584 ;
			LAYER M4 ;
			RECT 0.120 31.864 15.397 32.024 ;
			LAYER M4 ;
			RECT 0.120 33.304 15.397 33.464 ;
			LAYER M4 ;
			RECT 0.120 34.744 15.397 34.904 ;
			LAYER M4 ;
			RECT 0.120 36.184 15.397 36.344 ;
			LAYER M4 ;
			RECT 0.120 37.624 15.397 37.784 ;
			LAYER M4 ;
			RECT 0.120 39.064 15.397 39.224 ;
			LAYER M4 ;
			RECT 0.120 40.504 15.397 40.664 ;
			LAYER M4 ;
			RECT 0.120 41.944 15.397 42.104 ;
			LAYER M4 ;
			RECT 0.120 43.384 15.397 43.544 ;
			LAYER M4 ;
			RECT 0.120 44.824 15.397 44.984 ;
			LAYER M4 ;
			RECT 0.120 46.264 15.397 46.424 ;
			LAYER M4 ;
			RECT 0.120 47.684 15.397 47.884 ;
			LAYER M4 ;
			RECT 0.120 48.620 15.397 48.820 ;
			LAYER M4 ;
			RECT 0.120 50.156 15.397 50.356 ;
			LAYER M4 ;
			RECT 0.120 51.692 15.397 51.892 ;
			LAYER M4 ;
			RECT 0.120 53.228 15.397 53.428 ;
			LAYER M4 ;
			RECT 0.120 54.764 15.397 54.964 ;
			LAYER M4 ;
			RECT 0.120 56.300 15.397 56.500 ;
			LAYER M4 ;
			RECT 0.120 57.836 15.397 58.036 ;
			LAYER M4 ;
			RECT 0.120 59.372 15.397 59.572 ;
			LAYER M4 ;
			RECT 0.120 60.908 15.397 61.108 ;
			LAYER M4 ;
			RECT 0.120 62.444 15.397 62.644 ;
			LAYER M4 ;
			RECT 0.120 63.980 15.397 64.180 ;
			LAYER M4 ;
			RECT 0.120 64.916 15.397 65.116 ;
			LAYER M4 ;
			RECT 0.120 66.376 15.397 66.536 ;
			LAYER M4 ;
			RECT 0.120 67.816 15.397 67.976 ;
			LAYER M4 ;
			RECT 0.120 69.256 15.397 69.416 ;
			LAYER M4 ;
			RECT 0.120 70.696 15.397 70.856 ;
			LAYER M4 ;
			RECT 0.120 72.136 15.397 72.296 ;
			LAYER M4 ;
			RECT 0.120 73.576 15.397 73.736 ;
			LAYER M4 ;
			RECT 0.120 75.016 15.397 75.176 ;
			LAYER M4 ;
			RECT 0.120 76.456 15.397 76.616 ;
			LAYER M4 ;
			RECT 0.120 77.896 15.397 78.056 ;
			LAYER M4 ;
			RECT 0.120 79.336 15.397 79.496 ;
			LAYER M4 ;
			RECT 0.120 80.776 15.397 80.936 ;
			LAYER M4 ;
			RECT 0.120 82.216 15.397 82.376 ;
			LAYER M4 ;
			RECT 0.120 83.656 15.397 83.816 ;
			LAYER M4 ;
			RECT 0.120 85.096 15.397 85.256 ;
			LAYER M4 ;
			RECT 0.120 86.536 15.397 86.696 ;
			LAYER M4 ;
			RECT 0.120 87.976 15.397 88.136 ;
			LAYER M4 ;
			RECT 0.120 89.416 15.397 89.576 ;
			LAYER M4 ;
			RECT 0.120 90.856 15.397 91.016 ;
			LAYER M4 ;
			RECT 0.120 92.296 15.397 92.456 ;
			LAYER M4 ;
			RECT 0.120 93.736 15.397 93.896 ;
			LAYER M4 ;
			RECT 0.120 95.176 15.397 95.336 ;
			LAYER M4 ;
			RECT 0.120 96.616 15.397 96.776 ;
			LAYER M4 ;
			RECT 0.120 98.056 15.397 98.216 ;
			LAYER M4 ;
			RECT 0.120 99.496 15.397 99.656 ;
			LAYER M4 ;
			RECT 0.120 100.936 15.397 101.096 ;
			LAYER M4 ;
			RECT 0.120 102.376 15.397 102.536 ;
			LAYER M4 ;
			RECT 0.120 103.816 15.397 103.976 ;
			LAYER M4 ;
			RECT 0.120 105.256 15.397 105.416 ;
			LAYER M4 ;
			RECT 0.120 106.696 15.397 106.856 ;
			LAYER M4 ;
			RECT 0.120 108.136 15.397 108.296 ;
			LAYER M4 ;
			RECT 0.120 109.576 15.397 109.736 ;
			LAYER M4 ;
			RECT 0.120 111.016 15.397 111.176 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 0.884 15.397 1.084 ;
			LAYER M4 ;
			RECT 0.120 2.324 15.397 2.524 ;
			LAYER M4 ;
			RECT 0.120 3.764 15.397 3.964 ;
			LAYER M4 ;
			RECT 0.120 5.204 15.397 5.404 ;
			LAYER M4 ;
			RECT 0.120 6.644 15.397 6.844 ;
			LAYER M4 ;
			RECT 0.120 8.084 15.397 8.284 ;
			LAYER M4 ;
			RECT 0.120 9.524 15.397 9.724 ;
			LAYER M4 ;
			RECT 0.120 10.964 15.397 11.164 ;
			LAYER M4 ;
			RECT 0.120 12.404 15.397 12.604 ;
			LAYER M4 ;
			RECT 0.120 13.844 15.397 14.044 ;
			LAYER M4 ;
			RECT 0.120 15.284 15.397 15.484 ;
			LAYER M4 ;
			RECT 0.120 16.724 15.397 16.924 ;
			LAYER M4 ;
			RECT 0.120 18.164 15.397 18.364 ;
			LAYER M4 ;
			RECT 0.120 19.604 15.397 19.804 ;
			LAYER M4 ;
			RECT 0.120 21.044 15.397 21.244 ;
			LAYER M4 ;
			RECT 0.120 22.484 15.397 22.684 ;
			LAYER M4 ;
			RECT 0.120 23.924 15.397 24.124 ;
			LAYER M4 ;
			RECT 0.120 25.364 15.397 25.564 ;
			LAYER M4 ;
			RECT 0.120 26.804 15.397 27.004 ;
			LAYER M4 ;
			RECT 0.120 28.244 15.397 28.444 ;
			LAYER M4 ;
			RECT 0.120 29.684 15.397 29.884 ;
			LAYER M4 ;
			RECT 0.120 31.124 15.397 31.324 ;
			LAYER M4 ;
			RECT 0.120 32.564 15.397 32.764 ;
			LAYER M4 ;
			RECT 0.120 34.004 15.397 34.204 ;
			LAYER M4 ;
			RECT 0.120 35.444 15.397 35.644 ;
			LAYER M4 ;
			RECT 0.120 36.884 15.397 37.084 ;
			LAYER M4 ;
			RECT 0.120 38.324 15.397 38.524 ;
			LAYER M4 ;
			RECT 0.120 39.764 15.397 39.964 ;
			LAYER M4 ;
			RECT 0.120 41.204 15.397 41.404 ;
			LAYER M4 ;
			RECT 0.120 42.644 15.397 42.844 ;
			LAYER M4 ;
			RECT 0.120 44.084 15.397 44.284 ;
			LAYER M4 ;
			RECT 0.120 45.524 15.397 45.724 ;
			LAYER M4 ;
			RECT 0.120 46.964 15.397 47.164 ;
			LAYER M4 ;
			RECT 0.120 49.388 15.397 49.588 ;
			LAYER M4 ;
			RECT 0.120 50.924 15.397 51.124 ;
			LAYER M4 ;
			RECT 0.120 52.460 15.397 52.660 ;
			LAYER M4 ;
			RECT 0.120 53.996 15.397 54.196 ;
			LAYER M4 ;
			RECT 0.120 55.532 15.397 55.732 ;
			LAYER M4 ;
			RECT 0.120 57.068 15.397 57.268 ;
			LAYER M4 ;
			RECT 0.120 58.604 15.397 58.804 ;
			LAYER M4 ;
			RECT 0.120 60.140 15.397 60.340 ;
			LAYER M4 ;
			RECT 0.120 61.676 15.397 61.876 ;
			LAYER M4 ;
			RECT 0.120 63.212 15.397 63.412 ;
			LAYER M4 ;
			RECT 0.120 65.636 15.397 65.836 ;
			LAYER M4 ;
			RECT 0.120 67.076 15.397 67.276 ;
			LAYER M4 ;
			RECT 0.120 68.516 15.397 68.716 ;
			LAYER M4 ;
			RECT 0.120 69.956 15.397 70.156 ;
			LAYER M4 ;
			RECT 0.120 71.396 15.397 71.596 ;
			LAYER M4 ;
			RECT 0.120 72.836 15.397 73.036 ;
			LAYER M4 ;
			RECT 0.120 74.276 15.397 74.476 ;
			LAYER M4 ;
			RECT 0.120 75.716 15.397 75.916 ;
			LAYER M4 ;
			RECT 0.120 77.156 15.397 77.356 ;
			LAYER M4 ;
			RECT 0.120 78.596 15.397 78.796 ;
			LAYER M4 ;
			RECT 0.120 80.036 15.397 80.236 ;
			LAYER M4 ;
			RECT 0.120 81.476 15.397 81.676 ;
			LAYER M4 ;
			RECT 0.120 82.916 15.397 83.116 ;
			LAYER M4 ;
			RECT 0.120 84.356 15.397 84.556 ;
			LAYER M4 ;
			RECT 0.120 85.796 15.397 85.996 ;
			LAYER M4 ;
			RECT 0.120 87.236 15.397 87.436 ;
			LAYER M4 ;
			RECT 0.120 88.676 15.397 88.876 ;
			LAYER M4 ;
			RECT 0.120 90.116 15.397 90.316 ;
			LAYER M4 ;
			RECT 0.120 91.556 15.397 91.756 ;
			LAYER M4 ;
			RECT 0.120 92.996 15.397 93.196 ;
			LAYER M4 ;
			RECT 0.120 94.436 15.397 94.636 ;
			LAYER M4 ;
			RECT 0.120 95.876 15.397 96.076 ;
			LAYER M4 ;
			RECT 0.120 97.316 15.397 97.516 ;
			LAYER M4 ;
			RECT 0.120 98.756 15.397 98.956 ;
			LAYER M4 ;
			RECT 0.120 100.196 15.397 100.396 ;
			LAYER M4 ;
			RECT 0.120 101.636 15.397 101.836 ;
			LAYER M4 ;
			RECT 0.120 103.076 15.397 103.276 ;
			LAYER M4 ;
			RECT 0.120 104.516 15.397 104.716 ;
			LAYER M4 ;
			RECT 0.120 105.956 15.397 106.156 ;
			LAYER M4 ;
			RECT 0.120 107.396 15.397 107.596 ;
			LAYER M4 ;
			RECT 0.120 108.836 15.397 109.036 ;
			LAYER M4 ;
			RECT 0.120 110.276 15.397 110.476 ;
			LAYER M4 ;
			RECT 0.120 111.716 15.397 111.916 ;
		END
	END VSS

	PIN WCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 48.038 15.517 48.118 ;
			LAYER M2 ;
			RECT 15.269 48.038 15.517 48.118 ;
			LAYER M3 ;
			RECT 15.269 48.038 15.517 48.118 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[0]

	PIN WCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 47.810 15.517 47.890 ;
			LAYER M2 ;
			RECT 15.269 47.810 15.517 47.890 ;
			LAYER M3 ;
			RECT 15.269 47.810 15.517 47.890 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.269 51.230 15.517 51.310 ;
			LAYER M2 ;
			RECT 15.269 51.230 15.517 51.310 ;
			LAYER M3 ;
			RECT 15.269 51.230 15.517 51.310 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0886 LAYER M1 ;
		ANTENNAMAXAREACAR 9.6368 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0833 LAYER M2 ;
		ANTENNAMAXAREACAR 13.2425 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4593 LAYER M3 ;
		ANTENNAMAXAREACAR 211.0720 LAYER M3 ;
	END WEB

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 15.517 112.800 ;
		LAYER M2 ;
		RECT 0.000 0.000 15.517 112.800 ;
		LAYER M3 ;
		RECT 0.000 0.000 15.517 112.800 ;
		LAYER M4 ;
		RECT 0.227 0.524 14.967 0.724 ;
		LAYER M4 ;
		RECT 0.227 1.358 14.537 1.518 ;
		LAYER M4 ;
		RECT 0.227 1.890 14.537 2.050 ;
		LAYER M4 ;
		RECT 0.227 2.798 14.537 2.958 ;
		LAYER M4 ;
		RECT 0.227 3.330 14.537 3.490 ;
		LAYER M4 ;
		RECT 0.227 4.238 14.537 4.398 ;
		LAYER M4 ;
		RECT 0.227 4.770 14.537 4.930 ;
		LAYER M4 ;
		RECT 0.227 5.678 14.537 5.838 ;
		LAYER M4 ;
		RECT 0.227 6.210 14.537 6.370 ;
		LAYER M4 ;
		RECT 0.227 7.118 14.537 7.278 ;
		LAYER M4 ;
		RECT 0.227 7.650 14.537 7.810 ;
		LAYER M4 ;
		RECT 0.227 8.558 14.537 8.718 ;
		LAYER M4 ;
		RECT 0.227 9.090 14.537 9.250 ;
		LAYER M4 ;
		RECT 0.227 9.998 14.537 10.158 ;
		LAYER M4 ;
		RECT 0.227 10.530 14.537 10.690 ;
		LAYER M4 ;
		RECT 0.227 11.438 14.537 11.598 ;
		LAYER M4 ;
		RECT 0.227 11.970 14.537 12.130 ;
		LAYER M4 ;
		RECT 0.227 12.878 14.537 13.038 ;
		LAYER M4 ;
		RECT 0.227 13.410 14.537 13.570 ;
		LAYER M4 ;
		RECT 0.227 14.318 14.537 14.478 ;
		LAYER M4 ;
		RECT 0.227 14.850 14.537 15.010 ;
		LAYER M4 ;
		RECT 0.227 15.758 14.537 15.918 ;
		LAYER M4 ;
		RECT 0.227 16.290 14.537 16.450 ;
		LAYER M4 ;
		RECT 0.227 17.198 14.537 17.358 ;
		LAYER M4 ;
		RECT 0.227 17.730 14.537 17.890 ;
		LAYER M4 ;
		RECT 0.227 18.638 14.537 18.798 ;
		LAYER M4 ;
		RECT 0.227 19.170 14.537 19.330 ;
		LAYER M4 ;
		RECT 0.227 20.078 14.537 20.238 ;
		LAYER M4 ;
		RECT 0.227 20.610 14.537 20.770 ;
		LAYER M4 ;
		RECT 0.227 21.518 14.537 21.678 ;
		LAYER M4 ;
		RECT 0.227 22.050 14.537 22.210 ;
		LAYER M4 ;
		RECT 0.227 22.958 14.537 23.118 ;
		LAYER M4 ;
		RECT 0.227 23.490 14.537 23.650 ;
		LAYER M4 ;
		RECT 0.227 24.398 14.537 24.558 ;
		LAYER M4 ;
		RECT 0.227 24.930 14.537 25.090 ;
		LAYER M4 ;
		RECT 0.227 25.838 14.537 25.998 ;
		LAYER M4 ;
		RECT 0.227 26.370 14.537 26.530 ;
		LAYER M4 ;
		RECT 0.227 27.278 14.537 27.438 ;
		LAYER M4 ;
		RECT 0.227 27.810 14.537 27.970 ;
		LAYER M4 ;
		RECT 0.227 28.718 14.537 28.878 ;
		LAYER M4 ;
		RECT 0.227 29.250 14.537 29.410 ;
		LAYER M4 ;
		RECT 0.227 30.158 14.537 30.318 ;
		LAYER M4 ;
		RECT 0.227 30.690 14.537 30.850 ;
		LAYER M4 ;
		RECT 0.227 31.598 14.537 31.758 ;
		LAYER M4 ;
		RECT 0.227 32.130 14.537 32.290 ;
		LAYER M4 ;
		RECT 0.227 33.038 14.537 33.198 ;
		LAYER M4 ;
		RECT 0.227 33.570 14.537 33.730 ;
		LAYER M4 ;
		RECT 0.227 34.478 14.537 34.638 ;
		LAYER M4 ;
		RECT 0.227 35.010 14.537 35.170 ;
		LAYER M4 ;
		RECT 0.227 35.918 14.537 36.078 ;
		LAYER M4 ;
		RECT 0.227 36.450 14.537 36.610 ;
		LAYER M4 ;
		RECT 0.227 37.358 14.537 37.518 ;
		LAYER M4 ;
		RECT 0.227 37.890 14.537 38.050 ;
		LAYER M4 ;
		RECT 0.227 38.798 14.537 38.958 ;
		LAYER M4 ;
		RECT 0.227 39.330 14.537 39.490 ;
		LAYER M4 ;
		RECT 0.227 40.238 14.537 40.398 ;
		LAYER M4 ;
		RECT 0.227 40.770 14.537 40.930 ;
		LAYER M4 ;
		RECT 0.227 41.678 14.537 41.838 ;
		LAYER M4 ;
		RECT 0.227 42.210 14.537 42.370 ;
		LAYER M4 ;
		RECT 0.227 43.118 14.537 43.278 ;
		LAYER M4 ;
		RECT 0.227 43.650 14.537 43.810 ;
		LAYER M4 ;
		RECT 0.227 44.558 14.537 44.718 ;
		LAYER M4 ;
		RECT 0.227 45.090 14.537 45.250 ;
		LAYER M4 ;
		RECT 0.227 45.998 14.537 46.158 ;
		LAYER M4 ;
		RECT 0.227 46.530 14.537 46.690 ;
		LAYER M4 ;
		RECT 0.227 47.324 14.537 47.524 ;
		LAYER M4 ;
		RECT 0.227 48.236 14.537 48.436 ;
		LAYER M4 ;
		RECT 0.227 49.004 14.537 49.204 ;
		LAYER M4 ;
		RECT 0.227 49.772 14.537 49.972 ;
		LAYER M4 ;
		RECT 0.227 50.540 14.537 50.740 ;
		LAYER M4 ;
		RECT 0.227 51.308 14.537 51.508 ;
		LAYER M4 ;
		RECT 0.227 52.076 14.537 52.276 ;
		LAYER M4 ;
		RECT 0.227 52.844 14.537 53.044 ;
		LAYER M4 ;
		RECT 0.227 53.612 14.537 53.812 ;
		LAYER M4 ;
		RECT 0.227 54.380 14.537 54.580 ;
		LAYER M4 ;
		RECT 0.227 55.148 14.537 55.348 ;
		LAYER M4 ;
		RECT 0.227 55.916 14.537 56.116 ;
		LAYER M4 ;
		RECT 0.227 56.684 14.537 56.884 ;
		LAYER M4 ;
		RECT 0.227 57.452 14.537 57.652 ;
		LAYER M4 ;
		RECT 0.227 58.220 14.537 58.420 ;
		LAYER M4 ;
		RECT 0.227 58.988 14.537 59.188 ;
		LAYER M4 ;
		RECT 0.227 59.756 14.537 59.956 ;
		LAYER M4 ;
		RECT 0.227 60.524 14.537 60.724 ;
		LAYER M4 ;
		RECT 0.227 61.292 14.537 61.492 ;
		LAYER M4 ;
		RECT 0.227 62.060 14.537 62.260 ;
		LAYER M4 ;
		RECT 0.227 62.828 14.537 63.028 ;
		LAYER M4 ;
		RECT 0.227 63.596 14.537 63.796 ;
		LAYER M4 ;
		RECT 0.227 64.364 14.537 64.564 ;
		LAYER M4 ;
		RECT 0.227 65.276 14.537 65.476 ;
		LAYER M4 ;
		RECT 0.227 66.110 14.537 66.270 ;
		LAYER M4 ;
		RECT 0.227 66.642 14.537 66.802 ;
		LAYER M4 ;
		RECT 0.227 67.550 14.537 67.710 ;
		LAYER M4 ;
		RECT 0.227 68.082 14.537 68.242 ;
		LAYER M4 ;
		RECT 0.227 68.990 14.537 69.150 ;
		LAYER M4 ;
		RECT 0.227 69.522 14.537 69.682 ;
		LAYER M4 ;
		RECT 0.227 70.430 14.537 70.590 ;
		LAYER M4 ;
		RECT 0.227 70.962 14.537 71.122 ;
		LAYER M4 ;
		RECT 0.227 71.870 14.537 72.030 ;
		LAYER M4 ;
		RECT 0.227 72.402 14.537 72.562 ;
		LAYER M4 ;
		RECT 0.227 73.310 14.537 73.470 ;
		LAYER M4 ;
		RECT 0.227 73.842 14.537 74.002 ;
		LAYER M4 ;
		RECT 0.227 74.750 14.537 74.910 ;
		LAYER M4 ;
		RECT 0.227 75.282 14.537 75.442 ;
		LAYER M4 ;
		RECT 0.227 76.190 14.537 76.350 ;
		LAYER M4 ;
		RECT 0.227 76.722 14.537 76.882 ;
		LAYER M4 ;
		RECT 0.227 77.630 14.537 77.790 ;
		LAYER M4 ;
		RECT 0.227 78.162 14.537 78.322 ;
		LAYER M4 ;
		RECT 0.227 79.070 14.537 79.230 ;
		LAYER M4 ;
		RECT 0.227 79.602 14.537 79.762 ;
		LAYER M4 ;
		RECT 0.227 80.510 14.537 80.670 ;
		LAYER M4 ;
		RECT 0.227 81.042 14.537 81.202 ;
		LAYER M4 ;
		RECT 0.227 81.950 14.537 82.110 ;
		LAYER M4 ;
		RECT 0.227 82.482 14.537 82.642 ;
		LAYER M4 ;
		RECT 0.227 83.390 14.537 83.550 ;
		LAYER M4 ;
		RECT 0.227 83.922 14.537 84.082 ;
		LAYER M4 ;
		RECT 0.227 84.830 14.537 84.990 ;
		LAYER M4 ;
		RECT 0.227 85.362 14.537 85.522 ;
		LAYER M4 ;
		RECT 0.227 86.270 14.537 86.430 ;
		LAYER M4 ;
		RECT 0.227 86.802 14.537 86.962 ;
		LAYER M4 ;
		RECT 0.227 87.710 14.537 87.870 ;
		LAYER M4 ;
		RECT 0.227 88.242 14.537 88.402 ;
		LAYER M4 ;
		RECT 0.227 89.150 14.537 89.310 ;
		LAYER M4 ;
		RECT 0.227 89.682 14.537 89.842 ;
		LAYER M4 ;
		RECT 0.227 90.590 14.537 90.750 ;
		LAYER M4 ;
		RECT 0.227 91.122 14.537 91.282 ;
		LAYER M4 ;
		RECT 0.227 92.030 14.537 92.190 ;
		LAYER M4 ;
		RECT 0.227 92.562 14.537 92.722 ;
		LAYER M4 ;
		RECT 0.227 93.470 14.537 93.630 ;
		LAYER M4 ;
		RECT 0.227 94.002 14.537 94.162 ;
		LAYER M4 ;
		RECT 0.227 94.910 14.537 95.070 ;
		LAYER M4 ;
		RECT 0.227 95.442 14.537 95.602 ;
		LAYER M4 ;
		RECT 0.227 96.350 14.537 96.510 ;
		LAYER M4 ;
		RECT 0.227 96.882 14.537 97.042 ;
		LAYER M4 ;
		RECT 0.227 97.790 14.537 97.950 ;
		LAYER M4 ;
		RECT 0.227 98.322 14.537 98.482 ;
		LAYER M4 ;
		RECT 0.227 99.230 14.537 99.390 ;
		LAYER M4 ;
		RECT 0.227 99.762 14.537 99.922 ;
		LAYER M4 ;
		RECT 0.227 100.670 14.537 100.830 ;
		LAYER M4 ;
		RECT 0.227 101.202 14.537 101.362 ;
		LAYER M4 ;
		RECT 0.227 102.110 14.537 102.270 ;
		LAYER M4 ;
		RECT 0.227 102.642 14.537 102.802 ;
		LAYER M4 ;
		RECT 0.227 103.550 14.537 103.710 ;
		LAYER M4 ;
		RECT 0.227 104.082 14.537 104.242 ;
		LAYER M4 ;
		RECT 0.227 104.990 14.537 105.150 ;
		LAYER M4 ;
		RECT 0.227 105.522 14.537 105.682 ;
		LAYER M4 ;
		RECT 0.227 106.430 14.537 106.590 ;
		LAYER M4 ;
		RECT 0.227 106.962 14.537 107.122 ;
		LAYER M4 ;
		RECT 0.227 107.870 14.537 108.030 ;
		LAYER M4 ;
		RECT 0.227 108.402 14.537 108.562 ;
		LAYER M4 ;
		RECT 0.227 109.310 14.537 109.470 ;
		LAYER M4 ;
		RECT 0.227 109.842 14.537 110.002 ;
		LAYER M4 ;
		RECT 0.227 110.750 14.537 110.910 ;
		LAYER M4 ;
		RECT 0.227 111.282 14.537 111.442 ;
		LAYER M4 ;
		RECT 0.227 112.076 14.967 112.276 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 15.517 112.800 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 15.517 112.800 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 15.517 112.800 ;
	END
END TS6N16FFCLLSVTA32X32M4FW

END LIBRARY
