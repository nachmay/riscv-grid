**** Created by MC2: Version 2013.12.00.f on 2025/06/18, 12:59:41 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  TS16FF2PRF
* Top Cell Name: all_leafcells
* View Name:     schematic
* Netlisted on:  Sep 30 16:22:09 2015
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM


*.PIN vss

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_svt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nand2_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_svt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_inv_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_svt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nor2_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WCTD VDD VDDI VSS TSMC_1 TSMC_2 TSMC_3 TSMC_4 
XI76 TSMC_5 TSMC_6 VSS VSS VDDI VDD TSMC_3 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI79 TSMC_7 TSMC_8 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI66 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_2 TSMC_11 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_7 TSMC_12 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_14 TSMC_7 VSS VSS VDDI VDD TSMC_6 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_1 TSMC_15 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_9 TSMC_16 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_17 TSMC_11 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_16 TSMC_15 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI145 VSS VSS TSMC_4 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_18 TSMC_5 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_5 TSMC_19 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_5 TSMC_20 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI143 VSS VSS TSMC_21 TSMC_22 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI159 VSS VSS TSMC_13 TSMC_23 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_22 TSMC_17 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_24 TSMC_25 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI89 VSS VSS TSMC_10 TSMC_12 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI160 VSS VSS TSMC_13 TSMC_24 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI144 VSS VSS TSMC_25 TSMC_21 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW10V20_nor2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WRTRKEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WRTRKEN TSMC_1 VDD VDDI VSS TSMC_2 TSMC_3 TSMC_4 
XI19<0> TSMC_2 TSMC_5 VSS VSS VDDI VDD TSMC_1 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI19<1> TSMC_2 TSMC_5 VSS VSS VDDI VDD TSMC_1 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI14 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_5 
+ S6ALLSVTFW10V20_nor2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_W1TRKWR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_W1TRKWR TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS TSMC_4 
+ TSMC_5 
XXwctd VDD VDDI VSS TSMC_1 TSMC_2 TSMC_6 TSMC_4 S6ALLSVTFW10V20_RF_WCTD 
XXrdtrken TSMC_3 VDD VDDI VSS TSMC_6 TSMC_4 TSMC_5 
+ S6ALLSVTFW10V20_RF_WRTRKEN 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WREFMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WREFMUX TSMC_1 VDD VDDI VSS TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
MM10 TSMC_7 TSMC_1 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_4 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_4 TSMC_6 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM13 TSMC_8 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_3 TSMC_6 TSMC_9 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM12 TSMC_9 TSMC_1 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_3 TSMC_5 TSMC_4 VDD pch_svt_mac l=0.020u nfin=3 m=2 
MM9 TSMC_3 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM8 TSMC_4 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM0 TSMC_3 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_1 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_3 TSMC_10 TSMC_2 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM5 TSMC_4 TSMC_11 TSMC_2 VSS nch_svt_mac l=0.020u nfin=6 m=2 
XI21 TSMC_6 TSMC_7 TSMC_2 VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI19 TSMC_6 TSMC_1 TSMC_2 VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKGIOWR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TRKGIOWR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 
XXwrst TSMC_15 TSMC_16 TSMC_20 VDD VDDI VSS TSMC_17 TSMC_29 
+ S6ALLSVTFW10V20_RF_W1TRKWR 
XXwrefmux TSMC_11 VDD VDDI VSS VSS TSMC_12 TSMC_14 TSMC_30 TSMC_29 
+ S6ALLSVTFW10V20_RF_WREFMUX 
XI21 VSS VSS TSMC_19 TSMC_29 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_29 TSMC_30 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 p_nfin=7 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WMUX TSMC_1 TSMC_2 VDD VDDI VSS TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM0 TSMC_4 TSMC_8 TSMC_3 VSS nch_lvt_mac l=0.020u nfin=6 m=2 
MM2 TSMC_5 TSMC_9 TSMC_3 VSS nch_lvt_mac l=0.020u nfin=6 m=2 
MM13 TSMC_10 TSMC_1 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_4 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_4 TSMC_11 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_5 TSMC_11 TSMC_10 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM9 TSMC_4 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM4 TSMC_5 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM10 TSMC_4 TSMC_6 TSMC_5 VDD pch_svt_mac l=0.020u nfin=3 m=2 
MM6 TSMC_5 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM12 TSMC_12 TSMC_2 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI23 VSS VSS TSMC_7 TSMC_11 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI14 TSMC_11 TSMC_2 TSMC_3 VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI15 TSMC_11 TSMC_1 TSMC_3 VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRI_W3L2M1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TRI_W3L2M1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM4 TSMC_9 TSMC_7 TSMC_4 TSMC_5 pch_svt_mac l=0.020u nfin=3 m=1 
MM5 TSMC_8 TSMC_1 TSMC_9 TSMC_5 pch_svt_mac l=0.020u nfin=3 m=1 
MM6 TSMC_10 TSMC_6 TSMC_2 TSMC_3 nch_svt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_8 TSMC_1 TSMC_10 TSMC_3 nch_svt_mac l=0.020u nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRI_W2L2M1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TRI_W2L2M1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM4 TSMC_9 TSMC_7 TSMC_4 TSMC_5 pch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_8 TSMC_1 TSMC_9 TSMC_5 pch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_10 TSMC_6 TSMC_2 TSMC_3 nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_8 TSMC_1 TSMC_10 TSMC_3 nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DIN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_DIN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD 
+ VDDI VSS TSMC_7 
XI16 TSMC_8 VSS VSS VDDI VDD TSMC_4 TSMC_5 TSMC_9 
+ S6ALLSVTFW10V20_RF_TRI_W3L2M1 
XI90 TSMC_10 VSS VSS VDDI VDD TSMC_4 TSMC_5 TSMC_11 
+ S6ALLSVTFW10V20_RF_TRI_W3L2M1 
XI15 TSMC_12 TSMC_13 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_12 TSMC_14 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI63 VSS VSS TSMC_15 TSMC_12 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI59 VSS VSS TSMC_16 TSMC_14 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI61 VSS VSS TSMC_7 TSMC_17 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI83 VSS VSS TSMC_9 TSMC_3 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI92 VSS VSS TSMC_11 TSMC_2 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI99 VSS VSS TSMC_1 TSMC_16 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI62 VSS VSS TSMC_17 TSMC_15 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI60 VSS VSS TSMC_14 TSMC_13 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI94 TSMC_2 VSS VSS VDDI VDD TSMC_5 TSMC_4 TSMC_11 
+ S6ALLSVTFW10V20_RF_TRI_W2L2M1 
XI17 TSMC_3 VSS VSS VDDI VDD TSMC_5 TSMC_4 TSMC_9 
+ S6ALLSVTFW10V20_RF_TRI_W2L2M1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    TRI_M2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_TRI_M2 TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS TSMC_4 
MM4 TSMC_5 TSMC_1 VDDI VDD pch_lvt_mac l=0.020u nfin=4 m=1 
MM5 TSMC_4 TSMC_3 TSMC_5 VDD pch_lvt_mac l=0.020u nfin=4 m=1 
MM6 TSMC_6 TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=4 m=1 
MM3 TSMC_4 TSMC_2 TSMC_6 VSS nch_svt_mac l=0.020u nfin=4 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RMUX TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI VSS 
XI9 TSMC_1 TSMC_5 TSMC_4 VDD VDDI VSS TSMC_2 S6ALLSVTFW10V20_TRI_M2 
MM2 TSMC_1 TSMC_6 TSMC_7 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_7 TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_1 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=4 m=3 
MM5 TSMC_8 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_1 TSMC_6 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI1 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DOLATCH
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_DOLATCH TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 
MM2 TSMC_3 TSMC_4 VDD VDD pch_svt_mac l=0.020u nfin=3 m=1 
XI3 VSS VSS TSMC_3 TSMC_1 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI7 TSMC_2 VSS VSS VDDI VDD TSMC_5 TSMC_6 TSMC_3 
+ S6ALLSVTFW10V20_RF_TRI_W2L2M1 
XI5 TSMC_3 VSS VSS VDDI VDD TSMC_7 TSMC_8 TSMC_2 
+ S6ALLSVTFW10V20_RF_TRI_W2L2M1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DOUTM2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_DOUTM2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS TSMC_9 TSMC_10 
MM2 TSMC_11 TSMC_9 TSMC_12 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_12 TSMC_8 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
XXrmux_f TSMC_2 TSMC_13 TSMC_14 TSMC_15 TSMC_16 VDD VDDI VSS 
+ S6ALLSVTFW10V20_RF_RMUX 
XXrmux<0> TSMC_3 TSMC_13 TSMC_14 TSMC_17 TSMC_18 VDD VDDI VSS 
+ S6ALLSVTFW10V20_RF_RMUX 
XXqltch TSMC_5 TSMC_1 TSMC_13 TSMC_4 TSMC_19 TSMC_20 VDD VDDI VSS TSMC_9 
+ TSMC_10 S6ALLSVTFW10V20_RF_DOLATCH 
XI13 VSS VSS TSMC_20 TSMC_19 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_20 TSMC_21 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI6<1> VSS VSS TSMC_16 TSMC_15 VDD VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI6<0> VSS VSS TSMC_18 TSMC_17 VDD VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI7 VSS VSS TSMC_11 TSMC_22 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI18 VSS VSS TSMC_21 TSMC_14 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI20 TSMC_4 TSMC_11 VSS VSS VDD VDD TSMC_20 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI8<1> TSMC_6 TSMC_11 VSS VSS VDD VDD TSMC_16 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI8<0> TSMC_7 TSMC_11 VSS VSS VDD VDD TSMC_18 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
MM0 TSMC_11 TSMC_9 VDD VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_11 TSMC_8 VDD VDD pch_lvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DINM2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_DINM2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 
XXdltch TSMC_1 TSMC_2 TSMC_3 TSMC_16 TSMC_17 TSMC_4 VDD VDDI VSS TSMC_11 
+ S6ALLSVTFW10V20_RF_DIN 
XXwmux_f TSMC_2 TSMC_3 VDD VDDI VSS TSMC_5 TSMC_7 TSMC_9 TSMC_18 
+ TSMC_14 S6ALLSVTFW10V20_RF_WMUX 
XXwmux<0> TSMC_2 TSMC_3 VDD VDDI VSS TSMC_6 TSMC_8 TSMC_10 TSMC_18 
+ TSMC_15 S6ALLSVTFW10V20_RF_WMUX 
XI7 VSS VSS TSMC_19 TSMC_18 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 p_nfin=7 p_l=0.020u 
XI6 VSS VSS TSMC_13 TSMC_19 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI13 VSS VSS TSMC_12 TSMC_16 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI30 VSS VSS TSMC_16 TSMC_17 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_GIOM2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_GIOM2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDI VSS TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 
XXdout TSMC_2 TSMC_3 TSMC_4 TSMC_29 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS 
+ TSMC_14 TSMC_15 S6ALLSVTFW10V20_RF_DOUTM2 
XXdin TSMC_1 TSMC_5 TSMC_6 TSMC_12 VDD VDDI VSS TSMC_13 TSMC_13 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_27 TSMC_28 
+ S6ALLSVTFW10V20_RF_DINM2 
XI26 VSS VSS TSMC_7 TSMC_29 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_svt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nand3_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RLCTRL_DK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RLCTRL_DK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 VDD VDDI VSS TSMC_27 
MM12 TSMC_28 TSMC_29 TSMC_30 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM11 TSMC_30 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM7 TSMC_32 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM6 TSMC_33 TSMC_34 TSMC_32 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM5 TSMC_33 TSMC_35 TSMC_32 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM1 TSMC_36 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=8 m=16 
MM0 TSMC_36 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=8 m=16 
MM8 TSMC_28 TSMC_35 TSMC_30 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM13 TSMC_28 TSMC_31 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM4 TSMC_33 TSMC_31 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM3 TSMC_33 TSMC_35 TSMC_37 VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM2 TSMC_37 TSMC_34 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM10 TSMC_38 TSMC_29 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM9 TSMC_28 TSMC_35 TSMC_38 VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
XI96 TSMC_36 VSS TSMC_39 TSMC_18 VDD VDD 
+ S6ALLSVTFW10V20_inv_ulvt_mac_pcell n_totalM=16 n_nfin=6 n_l=0.020u 
+ p_totalM=16 p_nfin=6 p_l=0.020u 
XI100 VSS VSS TSMC_1 TSMC_40 VDDI VDD 
+ S6ALLSVTFW10V20_inv_ulvt_mac_pcell n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI107 VSS VSS TSMC_41 TSMC_5 VDD VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI91 VSS VSS TSMC_33 TSMC_42 VDD VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=5 n_nfin=7 n_l=0.020u p_totalM=5 p_nfin=6 p_l=0.020u 
XI92 TSMC_36 VSS TSMC_42 TSMC_19 VDD VDD 
+ S6ALLSVTFW10V20_inv_ulvt_mac_pcell n_totalM=16 n_nfin=6 n_l=0.020u 
+ p_totalM=16 p_nfin=6 p_l=0.020u 
XI106 VSS VSS TSMC_4 TSMC_41 VDD VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI98 VSS VSS TSMC_35 TSMC_23 VDDI VDD 
+ S6ALLSVTFW10V20_inv_ulvt_mac_pcell n_totalM=14 n_nfin=5 n_l=0.020u 
+ p_totalM=14 p_nfin=5 p_l=0.020u 
XI101 VSS VSS TSMC_40 TSMC_11 VDDI VDD 
+ S6ALLSVTFW10V20_inv_ulvt_mac_pcell n_totalM=10 n_nfin=7 n_l=0.020u 
+ p_totalM=10 p_nfin=8 p_l=0.020u 
XI93_Lg16 TSMC_21 TSMC_22 TSMC_27 VSS VSS VDD VDD TSMC_35 
+ S6ALLSVTFW10V20_nand3_ulvt_mac_pcell n_totalM=4 n_nfin=7 n_l=0.020u 
+ p_totalM=4 p_nfin=2 p_l=0.020u 
XI95 TSMC_25 TSMC_26 VSS VSS VDDI VDD TSMC_34 
+ S6ALLSVTFW10V20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI103 TSMC_28 TSMC_24 VSS VSS VDD VDD TSMC_39 
+ S6ALLSVTFW10V20_nor2_ulvt_mac_pcell n_totalM=6 n_nfin=6 n_l=0.020u p_totalM=6 
+ p_nfin=7 p_l=0.020u 
XI102 TSMC_4 TSMC_4 VSS VSS VDD VDD TSMC_31 
+ S6ALLSVTFW10V20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI99 TSMC_2 TSMC_3 VSS VSS VDDI VDD TSMC_29 
+ S6ALLSVTFW10V20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WLCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WLCTRL VDD VDDI VSS TSMC_1 TSMC_2 TSMC_3 TSMC_4 
XI27 TSMC_1 TSMC_2 TSMC_4 VSS VSS VDD VDD TSMC_5 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=4 n_nfin=7 n_l=0.020u p_totalM=4 
+ p_nfin=2 p_l=0.020u 
XI28 VSS VSS TSMC_5 TSMC_3 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=14 n_nfin=5 n_l=0.020u p_totalM=14 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LCTRL_DK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_LCTRL_DK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
MM6 TSMC_71 TSMC_46 VDD VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM4 VDDI TSMC_46 VDDI VDD pch_ulvt_mac l=0.020u nfin=8 m=2 
MM5 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=12 m=16 
MM1 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=5 m=16 
MM0 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=9 m=32 
MM2 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=10 m=16 
XXrlctrl TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_17 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_25 TSMC_27 TSMC_28 TSMC_45 TSMC_48 TSMC_49 VDD 
+ VDDI VSS TSMC_69 S6ALLSVTFW10V20_RF_RLCTRL_DK 
XXwlctrl VDD VDDI VSS TSMC_50 TSMC_51 TSMC_52 TSMC_70 
+ S6ALLSVTFW10V20_RF_WLCTRL 
XI51 VSS VSS TSMC_73 TSMC_72 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI52 TSMC_24 TSMC_4 VSS VSS VDD VDD TSMC_73 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
MM3 VSS TSMC_46 VSS VSS nch_ulvt_mac l=0.020u nfin=7 m=2 
MM7 TSMC_46 TSMC_71 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_LCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
XI152 TSMC_15 TSMC_24 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=2 n_nfin=12 n_l=0.020u p_totalM=2 
+ p_nfin=12 p_l=0.020u 
XI49<1> VSS VSS TSMC_18 TSMC_12 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI49<0> VSS VSS TSMC_19 TSMC_13 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
Xlctrl TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ S6ALLSVTFW10V20_RF_LCTRL_DK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_XDECCAP
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_XDECCAP TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 
MM0_LVT TSMC_12 TSMC_6 VSS VSS nch_lvt_mac l=0.020u nfin=5 m=1 
MM196_LVT TSMC_13 TSMC_12 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM197_LVT TSMC_14 TSMC_12 TSMC_13 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM194_LVT TSMC_12 TSMC_15 VSS VSS nch_lvt_mac l=0.020u nfin=5 m=1 
MM4 TSMC_10 TSMC_16 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MMWLDRPCHWTK TSMC_10 TSMC_16 VDDI VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM195_LVT TSMC_14 TSMC_12 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=2 
MM198_LVT TSMC_17 TSMC_15 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM193_LVT TSMC_12 TSMC_6 TSMC_17 VDD pch_lvt_mac l=0.020u nfin=2 m=1 
XI78 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=6 n_l=0.020u p_totalM=2 p_nfin=6 p_l=0.020u 
XI75 VSS VSS TSMC_9 TSMC_18 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI79 VSS VSS TSMC_3 TSMC_4 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI72_LVT VSS VSS TSMC_11 TSMC_15 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI73_LVT VSS VSS TSMC_14 TSMC_19 VDDI VDD 
+ S6ALLSVTFW10V20_inv_lvt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI77 VSS VSS TSMC_2 TSMC_20 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI76 VSS VSS TSMC_18 TSMC_21 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI81_LVT TSMC_10 TSMC_19 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=8 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI82 TSMC_20 TSMC_21 VSS VSS VDD VDD TSMC_16 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=12 n_l=0.020u 
+ p_totalM=1 p_nfin=10 p_l=0.020u 
XI80_LVT TSMC_10 TSMC_19 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=6 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TRKCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 VDD VDDI VSS TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 
MM4 TSMC_37 TSMC_56 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
XI76 VSS VSS TSMC_57 TSMC_58 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI75 VSS VSS TSMC_12 TSMC_57 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI78 TSMC_13 TSMC_14 VSS VSS VDD VDD TSMC_56 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=12 n_l=0.020u 
+ p_totalM=1 p_nfin=6 p_l=0.020u 
XI79 TSMC_58 TSMC_14 VSS VSS VDDI VDD TSMC_59 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=7 p_l=0.020u 
MMWLDRPCHRTK TSMC_37 TSMC_56 VDDI VDD pch_svt_mac l=0.020u nfin=11 m=4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WXDEC TSMC_1 TSMC_2 TSMC_3 VDD VDDI TSMC_4 VSS 
+ TSMC_5 TSMC_6 
MM3 TSMC_1 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM2 TSMC_7 TSMC_8 TSMC_1 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM4 TSMC_5 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MMWLDRPCH TSMC_5 TSMC_7 TSMC_4 VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MM0 TSMC_7 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
XI58<1> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI58<0> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDECX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WXDECX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XI64<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XIXDEC<3> TSMC_16 TSMC_2 TSMC_3 VDD VDDI TSMC_7 VSS TSMC_8 TSMC_15 
+ S6ALLSVTFW10V20_RF_WXDEC 
XIXDEC<1> TSMC_16 TSMC_2 TSMC_5 VDD VDDI TSMC_7 VSS TSMC_10 TSMC_15 
+ S6ALLSVTFW10V20_RF_WXDEC 
XIXDEC<0> TSMC_17 TSMC_1 TSMC_6 VDD VDDI TSMC_7 VSS TSMC_11 TSMC_14 
+ S6ALLSVTFW10V20_RF_WXDEC 
XIXDEC<2> TSMC_17 TSMC_1 TSMC_4 VDD VDDI TSMC_7 VSS TSMC_9 TSMC_14 
+ S6ALLSVTFW10V20_RF_WXDEC 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDECX4_LR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WXDECX4_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD VDDI TSMC_7 VSS 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ S6ALLSVTFW10V20_RF_WXDECX4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RXDEC TSMC_1 TSMC_2 TSMC_3 VDD VDDI TSMC_4 VSS 
+ TSMC_5 TSMC_6 
MM1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MMWLDRPCH TSMC_5 TSMC_7 TSMC_4 VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM0 TSMC_7 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MM4 TSMC_5 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MM2 TSMC_7 TSMC_8 TSMC_1 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM3 TSMC_1 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=6 m=2 
XI58<1> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI58<0> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDECX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RXDECX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC<1> TSMC_14 TSMC_2 TSMC_5 VDD VDDI TSMC_7 VSS TSMC_10 TSMC_15 
+ S6ALLSVTFW10V20_RF_RXDEC 
XIXDEC<3> TSMC_14 TSMC_2 TSMC_3 VDD VDDI TSMC_7 VSS TSMC_8 TSMC_15 
+ S6ALLSVTFW10V20_RF_RXDEC 
XIXDEC<2> TSMC_16 TSMC_1 TSMC_4 VDD VDDI TSMC_7 VSS TSMC_9 TSMC_17 
+ S6ALLSVTFW10V20_RF_RXDEC 
XIXDEC<0> TSMC_16 TSMC_1 TSMC_6 VDD VDDI TSMC_7 VSS TSMC_11 TSMC_17 
+ S6ALLSVTFW10V20_RF_RXDEC 
XI64<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDECX4_LR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RXDECX4_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD VDDI TSMC_7 VSS 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ S6ALLSVTFW10V20_RF_RXDECX4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_XDEC4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_XDEC4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 VDD VDDI TSMC_42 VSS 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
XXwdec TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 VDD VDDI TSMC_42 VSS 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_69 TSMC_70 
+ S6ALLSVTFW10V20_RF_WXDECX4_LR 
XXrdec TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 VDD VDDI TSMC_42 VSS 
+ TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_67 TSMC_68 
+ S6ALLSVTFW10V20_RF_RXDECX4_LR 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TIELGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TIELGEN TSMC_1 TSMC_2 VDD VSS 
MM5 TSMC_1 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_3 TSMC_4 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_2 TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=3 m=2 
MM2 TSMC_3 TSMC_5 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_2 TSMC_6 VSS VSS nch_svt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_3 TSMC_5 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI0 VSS VSS TSMC_5 TSMC_4 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI1 VSS VSS TSMC_4 TSMC_6 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PUDELAY
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_PUDELAY TSMC_1 TSMC_2 TSMC_3 VDD VSS 
XI3 VSS VSS TSMC_4 TSMC_2 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI149 TSMC_1 TSMC_3 VSS VSS VDD VDD TSMC_4 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DEC2TO4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_DEC2TO4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS 
XI26 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI27 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI28 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI33 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI34 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI37 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI31 VSS VSS TSMC_10 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI35 VSS VSS TSMC_11 TSMC_6 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI39 VSS VSS TSMC_12 TSMC_5 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI29 VSS VSS TSMC_9 TSMC_8 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_YDEC3TO8L
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_YDEC3TO8L TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
XI32 TSMC_3 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI42 TSMC_6 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI38 TSMC_6 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI43 TSMC_3 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI39 TSMC_3 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_19 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI35 TSMC_6 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_3 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_6 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 VSS VSS TSMC_17 TSMC_23 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI82 VSS VSS TSMC_24 TSMC_12 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI15 VSS VSS TSMC_25 TSMC_14 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI85 VSS VSS TSMC_26 TSMC_9 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI3 VSS VSS TSMC_22 TSMC_25 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI94 VSS VSS TSMC_18 TSMC_27 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI93 VSS VSS TSMC_16 TSMC_28 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI81 VSS VSS TSMC_29 TSMC_13 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI87 VSS VSS TSMC_27 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI92 VSS VSS TSMC_19 TSMC_26 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI90 VSS VSS TSMC_21 TSMC_30 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI83 VSS VSS TSMC_30 TSMC_11 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI84 VSS VSS TSMC_23 TSMC_10 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI89 VSS VSS TSMC_20 TSMC_24 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI88 VSS VSS TSMC_15 TSMC_29 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI86 VSS VSS TSMC_28 TSMC_8 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DECPDA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_DECPDA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS 
XI58 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI60 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI59 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI61 VSS VSS TSMC_9 TSMC_13 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI64 VSS VSS TSMC_11 TSMC_14 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI66 VSS VSS TSMC_15 TSMC_5 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI62 VSS VSS TSMC_13 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI63 VSS VSS TSMC_14 TSMC_6 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI65 VSS VSS TSMC_10 TSMC_15 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI35 VSS VSS TSMC_16 TSMC_8 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI42 VSS VSS TSMC_12 TSMC_16 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RPREDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RPREDEC TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI VSS TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 
XXpb TSMC_5 TSMC_6 TSMC_13 TSMC_14 TSMC_27 TSMC_28 TSMC_29 TSMC_30 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DEC2TO4 
XXpd TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DEC2TO4 
XXpc TSMC_3 TSMC_4 TSMC_11 TSMC_12 TSMC_31 TSMC_32 TSMC_33 TSMC_34 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DEC2TO4 
XXya TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 VDD VDDI VSS TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ S6ALLSVTFW10V20_RF_YDEC3TO8L 
XXpa TSMC_7 TSMC_8 TSMC_15 TSMC_16 TSMC_23 TSMC_24 TSMC_25 TSMC_26 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DECPDA 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RPRCHBUF
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RPRCHBUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_1 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI43 VSS VSS TSMC_3 TSMC_7 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=6 n_l=0.020u p_totalM=3 p_nfin=4 p_l=0.020u 
XI42 VSS VSS TSMC_1 TSMC_2 TSMC_6 VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI2 VSS VSS TSMC_7 TSMC_4 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=13 n_nfin=5 n_l=0.020u p_totalM=13 p_nfin=9 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RCLKGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RCLKGEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS 
XI53 TSMC_11 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW10V20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=8 p_l=0.016u 
XI25 TSMC_13 TSMC_2 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
XI73 VSS VSS TSMC_9 TSMC_15 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI5 VSS VSS TSMC_13 TSMC_16 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI6 VSS VSS TSMC_13 TSMC_3 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=9 n_nfin=5 n_l=0.016u p_totalM=9 p_nfin=5 p_l=0.016u 
XI40 VSS VSS TSMC_12 TSMC_17 VDDI VDD 
+ S6ALLSVTFW10V20_inv_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI2 VSS VSS TSMC_18 TSMC_19 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI29 VSS VSS TSMC_2 TSMC_20 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI19 VSS VSS TSMC_1 TSMC_2 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI79 VSS VSS TSMC_7 TSMC_6 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=2 n_nfin=5 n_l=0.016u p_totalM=2 p_nfin=5 p_l=0.016u 
XI17 VSS VSS TSMC_15 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=2 n_nfin=8 n_l=0.016u p_totalM=2 p_nfin=8 p_l=0.016u 
MM1 TSMC_21 TSMC_22 VDD VDD pch_ulvt_mac l=0.016u nfin=8 m=3 
MM3 TSMC_13 TSMC_4 TSMC_21 VDD pch_ulvt_mac l=0.016u nfin=8 m=3 
MM9 TSMC_18 TSMC_8 TSMC_23 VDD pch_ulvt_mac l=0.016u nfin=6 m=1 
MM5 TSMC_23 TSMC_20 VDDI VDD pch_ulvt_mac l=0.016u nfin=6 m=1 
MM13 TSMC_24 TSMC_12 VDD VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM6 TSMC_18 TSMC_19 TSMC_25 VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM12 TSMC_13 TSMC_16 TSMC_24 VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM10 TSMC_25 TSMC_14 VDDI VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM0 TSMC_16 TSMC_8 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=2 
MM8 TSMC_13 TSMC_12 VSS VSS nch_ulvt_mac l=0.016u nfin=5 m=6 
MM4 TSMC_26 TSMC_20 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM11 TSMC_18 TSMC_8 VSS VSS nch_ulvt_mac l=0.016u nfin=4 m=1 
MM2 TSMC_18 TSMC_14 VSS VSS nch_ulvt_mac l=0.016u nfin=4 m=1 
MM15 TSMC_27 TSMC_16 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM7 TSMC_18 TSMC_19 TSMC_26 VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM14 TSMC_13 TSMC_16 TSMC_27 VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
XI71 TSMC_13 TSMC_28 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nand2_ulvt_mac_pcell n_totalM=2 n_nfin=3 n_l=0.016u 
+ p_totalM=2 p_nfin=3 p_l=0.016u 
XI75 TSMC_5 TSMC_20 VSS VSS VDD VDD TSMC_28 
+ S6ALLSVTFW10V20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u 
+ p_totalM=1 p_nfin=2 p_l=0.016u 
XI56 TSMC_18 TSMC_5 VSS VSS VDD VDD TSMC_11 
+ S6ALLSVTFW10V20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u 
+ p_totalM=1 p_nfin=2 p_l=0.016u 
XI82 TSMC_29 TSMC_17 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW10V20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u 
+ p_totalM=1 p_nfin=3 p_l=0.016u 
XI8 TSMC_20 TSMC_10 VSS VSS VDDI VDD TSMC_29 
+ S6ALLSVTFW10V20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u 
+ p_totalM=1 p_nfin=2 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH_RA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_ILATCH_RA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_ulvt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_ulvt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW10V20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_ulvt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_ulvt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH_RA_Y
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_ILATCH_RA_Y TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_lvt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_lvt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW10V20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_lvt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_lvt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ADRLAT_RA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_ADRLAT_RA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 VDD VDDI VSS 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 
XXxlat<7> TSMC_25 TSMC_1 TSMC_2 TSMC_3 TSMC_11 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXxlat<6> TSMC_26 TSMC_1 TSMC_2 TSMC_4 TSMC_12 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXxlat<5> TSMC_27 TSMC_1 TSMC_2 TSMC_5 TSMC_13 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXxlat<4> TSMC_28 TSMC_1 TSMC_2 TSMC_6 TSMC_14 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXxlat<3> TSMC_29 TSMC_1 TSMC_2 TSMC_7 TSMC_15 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXxlat<2> TSMC_30 TSMC_1 TSMC_2 TSMC_8 TSMC_16 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXxlat<1> TSMC_31 TSMC_1 TSMC_2 TSMC_9 TSMC_17 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXxlat<0> TSMC_32 TSMC_1 TSMC_2 TSMC_10 TSMC_18 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA 
XXylat<2> TSMC_33 TSMC_1 TSMC_2 TSMC_19 TSMC_22 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA_Y 
XXylat<1> TSMC_34 TSMC_1 TSMC_2 TSMC_20 TSMC_23 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA_Y 
XXylat<0> TSMC_35 TSMC_1 TSMC_2 TSMC_21 TSMC_24 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH_RA_Y 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RENLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RENLAT TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
XI15 VSS VSS TSMC_5 TSMC_3 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI0 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI5 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
MM4 TSMC_8 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_9 TSMC_5 TSMC_8 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_10 TSMC_6 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_9 TSMC_2 TSMC_10 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_9 TSMC_5 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_11 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_9 TSMC_2 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_12 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI6 TSMC_4 TSMC_9 VSS VSS VDD VDD TSMC_5 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RTUNE
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RTUNE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDI VSS 
XXenlat TSMC_1 TSMC_10 TSMC_8 TSMC_9 VDD VDDI VSS 
+ S6ALLSVTFW10V20_RF_RENLAT 
XI12<2> VSS VSS TSMC_13 TSMC_5 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI12<1> VSS VSS TSMC_14 TSMC_6 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI12<0> VSS VSS TSMC_15 TSMC_7 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI13<2> VSS VSS TSMC_2 TSMC_13 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI13<1> VSS VSS TSMC_3 TSMC_14 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI13<0> VSS VSS TSMC_4 TSMC_15 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI7 VSS VSS TSMC_11 TSMC_12 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=5 n_l=0.020u p_totalM=4 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RGCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RGCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 VDD VDDI VSS TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
XXpredecs TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
+ TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 VDD VDDI VSS TSMC_58 
+ TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ S6ALLSVTFW10V20_RF_RPREDEC 
XXrprchb TSMC_38 TSMC_82 TSMC_83 TSMC_43 TSMC_46 VDD VDDI VSS 
+ S6ALLSVTFW10V20_RF_RPRCHBUF 
XXclkgen TSMC_1 TSMC_84 TSMC_40 TSMC_44 TSMC_85 TSMC_8 TSMC_9 TSMC_38 TSMC_83 
+ TSMC_45 VDD VDDI VSS S6ALLSVTFW10V20_RF_RCLKGEN 
XXadrlat TSMC_8 TSMC_9 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 VDD VDDI VSS 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 S6ALLSVTFW10V20_RF_ADRLAT_RA 
XXrtune TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_85 
+ TSMC_82 TSMC_39 TSMC_41 TSMC_42 VDD VDDI VSS S6ALLSVTFW10V20_RF_RTUNE 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DKCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_DKCTD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM2 VDDI TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=4 m=1 
MM1 VSS TSMC_5 VSS VSS nch_svt_mac l=0.020u nfin=4 m=1 
XI126 TSMC_4 TSMC_5 VSS VSS VDDI VDD TSMC_6 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI64 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_7 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI76 TSMC_8 TSMC_9 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI66 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_12 TSMC_6 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI179 TSMC_14 TSMC_6 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI178 TSMC_16 TSMC_6 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_1 TSMC_18 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_2 TSMC_19 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI156 TSMC_6 TSMC_10 VSS VSS VDDI VDD TSMC_3 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=6 n_nfin=10 n_l=0.020u 
+ p_totalM=6 p_nfin=5 p_l=0.020u 
XI89 VSS VSS TSMC_11 TSMC_12 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_7 TSMC_8 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_15 TSMC_20 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_21 TSMC_19 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_17 TSMC_22 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_20 TSMC_18 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_22 TSMC_9 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_13 TSMC_21 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WCLKGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WCLKGEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS TSMC_9 
MM11 TSMC_10 TSMC_11 TSMC_12 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM10 TSMC_12 TSMC_13 VDDI VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM13 TSMC_14 TSMC_15 VDD VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM2 TSMC_16 TSMC_17 VDDI VDD pch_svt_mac l=0.016u nfin=6 m=1 
MM3 TSMC_18 TSMC_3 TSMC_19 VDD pch_svt_mac l=0.016u nfin=8 m=3 
MM1 TSMC_19 TSMC_20 VDD VDD pch_svt_mac l=0.016u nfin=8 m=3 
MM0 TSMC_10 TSMC_7 TSMC_16 VDD pch_svt_mac l=0.016u nfin=6 m=1 
MM12 TSMC_18 TSMC_21 TSMC_14 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM15 TSMC_22 TSMC_21 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM7 TSMC_10 TSMC_11 TSMC_23 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM14 TSMC_18 TSMC_21 TSMC_22 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM4 TSMC_23 TSMC_17 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM9 TSMC_21 TSMC_7 VSS VSS nch_svt_mac l=0.016u nfin=2 m=2 
MM8 TSMC_18 TSMC_15 VSS VSS nch_svt_mac l=0.016u nfin=5 m=6 
MM5 TSMC_10 TSMC_7 VSS VSS nch_svt_mac l=0.016u nfin=4 m=1 
MM6 TSMC_10 TSMC_13 VSS VSS nch_svt_mac l=0.016u nfin=4 m=1 
XI61 VSS VSS TSMC_24 TSMC_9 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=5 n_l=0.016u p_totalM=6 p_nfin=5 p_l=0.016u 
XI48 VSS VSS TSMC_18 TSMC_6 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=8 n_l=0.016u p_totalM=3 p_nfin=9 p_l=0.016u 
XI45 VSS VSS TSMC_18 TSMC_25 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI28 VSS VSS TSMC_26 TSMC_24 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=8 n_l=0.016u p_totalM=1 p_nfin=8 p_l=0.016u 
XI17 VSS VSS TSMC_6 TSMC_5 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=8 n_l=0.016u p_totalM=1 p_nfin=8 p_l=0.016u 
XI44 VSS VSS TSMC_25 TSMC_27 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.016u p_totalM=2 p_nfin=4 p_l=0.016u 
XI5 VSS VSS TSMC_18 TSMC_21 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI29 VSS VSS TSMC_18 TSMC_26 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI6 VSS VSS TSMC_27 TSMC_2 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=5 n_l=0.016u p_totalM=6 p_nfin=5 p_l=0.016u 
XI26 VSS VSS TSMC_24 TSMC_9 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.016u p_totalM=4 p_nfin=8 p_l=0.016u 
XI2 VSS VSS TSMC_10 TSMC_11 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI1 VSS VSS TSMC_28 TSMC_17 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI0 VSS VSS TSMC_1 TSMC_28 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI40 VSS VSS TSMC_15 TSMC_29 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI8 TSMC_17 TSMC_8 VSS VSS VDDI VDD TSMC_30 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI37 TSMC_30 TSMC_29 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
XI52 TSMC_10 TSMC_4 VSS VSS VDD VDD TSMC_31 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI53 TSMC_31 TSMC_28 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=8 p_l=0.016u 
XI50 TSMC_18 TSMC_28 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_YDEC3TO8
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_YDEC3TO8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
XI32 TSMC_3 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI35 TSMC_6 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_3 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI38 TSMC_6 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI39 TSMC_3 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_19 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI42 TSMC_6 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI43 TSMC_3 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_6 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI33 VSS VSS TSMC_15 TSMC_13 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI34 VSS VSS TSMC_16 TSMC_12 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI37 VSS VSS TSMC_17 TSMC_11 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI40 VSS VSS TSMC_18 TSMC_10 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI41 VSS VSS TSMC_19 TSMC_9 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI44 VSS VSS TSMC_20 TSMC_8 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI29 VSS VSS TSMC_22 TSMC_14 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI45 VSS VSS TSMC_21 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WPREDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WPREDEC TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI VSS TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 
XXya TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 VDD VDDI VSS TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ S6ALLSVTFW10V20_RF_YDEC3TO8 
XXpb TSMC_5 TSMC_6 TSMC_13 TSMC_14 TSMC_27 TSMC_28 TSMC_29 TSMC_30 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DEC2TO4 
XXpd TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DEC2TO4 
XXpc TSMC_3 TSMC_4 TSMC_11 TSMC_12 TSMC_31 TSMC_32 TSMC_33 TSMC_34 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DEC2TO4 
XXpa TSMC_7 TSMC_8 TSMC_15 TSMC_16 TSMC_23 TSMC_24 TSMC_25 TSMC_26 VDD VDDI 
+ VSS S6ALLSVTFW10V20_RF_DECPDA 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ENLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_ENLAT TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS 
XI0 VSS VSS TSMC_1 TSMC_4 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI6 VSS VSS TSMC_5 TSMC_6 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI5 VSS VSS TSMC_4 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI4 VSS VSS TSMC_6 TSMC_3 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
MM5 TSMC_5 TSMC_6 TSMC_8 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_8 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_5 TSMC_2 TSMC_9 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_9 TSMC_4 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_5 TSMC_6 TSMC_10 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_10 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_5 TSMC_2 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_11 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WTUNE
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WTUNE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS TSMC_9 TSMC_10 TSMC_11 
XXenlat TSMC_1 TSMC_9 TSMC_8 VDD VDDI VSS S6ALLSVTFW10V20_RF_ENLAT 
XI15 VSS VSS TSMC_10 TSMC_11 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=7 n_l=0.020u p_totalM=3 p_nfin=7 p_l=0.020u 
XI9<2> VSS VSS TSMC_2 TSMC_12 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI9<1> VSS VSS TSMC_3 TSMC_13 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI9<0> VSS VSS TSMC_4 TSMC_14 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI8<2> VSS VSS TSMC_12 TSMC_5 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI8<1> VSS VSS TSMC_13 TSMC_6 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI8<0> VSS VSS TSMC_14 TSMC_7 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WPRCHBUF
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WPRCHBUF TSMC_1 TSMC_2 VDD VDDI VSS TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
XI18 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=7 p_l=0.020u 
XI17<7> TSMC_8 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<6> TSMC_9 TSMC_1 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<5> TSMC_10 TSMC_1 VSS VSS VDDI VDD TSMC_23 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<4> TSMC_11 TSMC_1 VSS VSS VDDI VDD TSMC_24 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<3> TSMC_4 TSMC_1 VSS VSS VDDI VDD TSMC_25 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<2> TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_26 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<1> TSMC_6 TSMC_1 VSS VSS VDDI VDD TSMC_27 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<0> TSMC_7 TSMC_1 VSS VSS VDDI VDD TSMC_28 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<7> TSMC_8 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<6> TSMC_9 TSMC_1 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<5> TSMC_10 TSMC_1 VSS VSS VDDI VDD TSMC_23 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<4> TSMC_11 TSMC_1 VSS VSS VDDI VDD TSMC_24 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<3> TSMC_4 TSMC_1 VSS VSS VDDI VDD TSMC_25 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<2> TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_26 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<1> TSMC_6 TSMC_1 VSS VSS VDDI VDD TSMC_27 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<0> TSMC_7 TSMC_1 VSS VSS VDDI VDD TSMC_28 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI7<7> VSS VSS TSMC_21 TSMC_12 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<6> VSS VSS TSMC_22 TSMC_13 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<5> VSS VSS TSMC_23 TSMC_14 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<4> VSS VSS TSMC_24 TSMC_15 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<3> VSS VSS TSMC_25 TSMC_16 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<2> VSS VSS TSMC_26 TSMC_17 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<1> VSS VSS TSMC_27 TSMC_18 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<0> VSS VSS TSMC_28 TSMC_19 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI2 VSS VSS TSMC_20 TSMC_3 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=9 n_l=16.0n p_totalM=6 p_nfin=9 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_ILATCH TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_svt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_svt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ADRLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_ADRLAT TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 VDD VDDI VSS 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 
XXylat<2> TSMC_33 TSMC_1 TSMC_2 TSMC_19 TSMC_22 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXylat<1> TSMC_34 TSMC_1 TSMC_2 TSMC_20 TSMC_23 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXylat<0> TSMC_35 TSMC_1 TSMC_2 TSMC_21 TSMC_24 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<7> TSMC_25 TSMC_1 TSMC_2 TSMC_3 TSMC_11 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<6> TSMC_26 TSMC_1 TSMC_2 TSMC_4 TSMC_12 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<5> TSMC_27 TSMC_1 TSMC_2 TSMC_5 TSMC_13 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<4> TSMC_28 TSMC_1 TSMC_2 TSMC_6 TSMC_14 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<3> TSMC_29 TSMC_1 TSMC_2 TSMC_7 TSMC_15 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<2> TSMC_30 TSMC_1 TSMC_2 TSMC_8 TSMC_16 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<1> TSMC_31 TSMC_1 TSMC_2 TSMC_9 TSMC_17 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
XXxlat<0> TSMC_32 TSMC_1 TSMC_2 TSMC_10 TSMC_18 VDD VDDI VSS 
+ S6ALLSVTFW10V20_ILATCH 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WGCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WGCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 VDD VDDI VSS TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 
XXclkgen TSMC_1 TSMC_33 TSMC_38 TSMC_62 TSMC_8 TSMC_9 TSMC_26 TSMC_31 VDD VDDI 
+ VSS TSMC_36 S6ALLSVTFW10V20_RF_WCLKGEN 
XXpredecs TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_10 TSMC_11 
+ TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 VDD VDDI VSS TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ S6ALLSVTFW10V20_RF_WPREDEC 
XXwtune TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_62 VDD VDDI VSS 
+ TSMC_32 TSMC_34 TSMC_35 S6ALLSVTFW10V20_RF_WTUNE 
XXwprchb TSMC_9 TSMC_26 VDD VDDI VSS TSMC_37 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 S6ALLSVTFW10V20_RF_WPRCHBUF 
XXadrlat TSMC_8 TSMC_9 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 VDD VDDI VSS 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 S6ALLSVTFW10V20_RF_ADRLAT 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_GCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_GCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 VDD VDDI VSS TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 
XXtiel TSMC_87 TSMC_88 VDD VSS S6ALLSVTFW10V20_RF_TIELGEN 
XXpudelay TSMC_27 TSMC_30 TSMC_86 VDD VSS S6ALLSVTFW10V20_RF_PUDELAY 
XXrctrl TSMC_1 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_20 
+ TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_29 TSMC_35 TSMC_36 TSMC_37 
+ TSMC_38 TSMC_71 TSMC_73 TSMC_89 TSMC_90 VDD VDDI VSS TSMC_75 TSMC_76 
+ TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 
+ TSMC_85 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 S6ALLSVTFW10V20_RF_RGCTRL 
XXdkctd TSMC_8 TSMC_9 TSMC_3 TSMC_13 TSMC_7 VDD VDDI VSS 
+ S6ALLSVTFW10V20_RF_DKCTD 
XXwctrl TSMC_2 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_29 TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_89 VDD VDDI VSS 
+ TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 
+ S6ALLSVTFW10V20_RF_WGCTRL 
MM1_header VDDI TSMC_28 VDD VDD pch_svt_mac l=0.020u nfin=7 m=24 
XI13 VSS VSS TSMC_28 TSMC_139 VDD VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI29 VSS VSS TSMC_88 TSMC_140 VDD VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=6 n_l=0.020u p_totalM=1 
+ p_nfin=6 p_l=0.020u 
XI3 VSS VSS TSMC_140 TSMC_141 VDD VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=2 n_nfin=6 n_l=0.020u p_totalM=2 
+ p_nfin=6 p_l=0.020u 
XI12 VSS VSS TSMC_139 TSMC_29 VDD VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=8 n_nfin=5 n_l=0.020u p_totalM=8 
+ p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PIN_GIO_MUX2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VSS 
XD5 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD4 VSS TSMC_2 ndio_mac nfin=2 l=200.0n m=1 
XD6 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD1 VSS TSMC_3 ndio_mac nfin=2 l=200.0n m=1 
XD2 VSS TSMC_4 ndio_mac nfin=2 l=200.0n m=1 
XD3 VSS TSMC_1 ndio_mac nfin=2 l=200.0n m=1 
XD7 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD8 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RCTD TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
XI79 TSMC_5 TSMC_6 VSS VSS VDDI VDD TSMC_7 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_2 TSMC_8 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_9 TSMC_6 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI76 TSMC_11 TSMC_10 VSS VSS VDDI VDD TSMC_4 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_12 TSMC_6 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI66 TSMC_2 TSMC_3 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_3 TSMC_15 VSS VSS VDDI VDD TSMC_5 
+ S6ALLSVTFW10V20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI149 VSS VSS TSMC_13 TSMC_16 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_11 TSMC_17 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI89 VSS VSS TSMC_14 TSMC_12 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_7 TSMC_18 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_19 TSMC_20 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_18 TSMC_8 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_21 TSMC_11 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_20 TSMC_15 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI145 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_11 TSMC_22 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI144 VSS VSS TSMC_23 TSMC_24 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI150 VSS VSS TSMC_13 TSMC_25 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_16 TSMC_23 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI143 VSS VSS TSMC_24 TSMC_19 VDDI VDD 
+ S6ALLSVTFW10V20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RDTRKEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_RDTRKEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS 
MM24 TSMC_11 TSMC_10 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM17 TSMC_4 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=4 m=4 
MM16 TSMC_4 TSMC_10 TSMC_12 VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM15 TSMC_12 TSMC_6 VSS VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM13 TSMC_3 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM8 TSMC_2 TSMC_10 TSMC_13 VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM2 TSMC_1 TSMC_14 TSMC_15 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM4 TSMC_15 TSMC_9 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM9 TSMC_16 TSMC_5 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM7 TSMC_13 TSMC_1 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM10 TSMC_3 TSMC_10 TSMC_16 VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM23 TSMC_2 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM3 VDDI TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM30 TSMC_10 TSMC_11 VDD VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM27 TSMC_2 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM20 TSMC_17 TSMC_6 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM19 TSMC_4 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=6 
MM18 TSMC_4 TSMC_11 TSMC_17 VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM14 TSMC_3 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM26 TSMC_3 TSMC_11 TSMC_18 VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM5 TSMC_19 TSMC_14 VDDI VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM0 TSMC_1 TSMC_14 TSMC_19 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM29 TSMC_2 TSMC_11 TSMC_20 VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM28 TSMC_20 TSMC_1 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM25 TSMC_18 TSMC_5 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM1 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.016u nfin=5 m=2 
XI33 TSMC_7 TSMC_2 TSMC_9 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW10V20_nand3_svt_mac_pcell n_totalM=2 n_nfin=6 n_l=0.016u p_totalM=2 
+ p_nfin=3 p_l=0.016u 
XI1 VSS VSS TSMC_1 TSMC_14 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKGIORD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TRKGIORD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 VDD VDDI VSS TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
XXrctd TSMC_4 TSMC_8 TSMC_9 TSMC_34 VDD VDDI VSS 
+ S6ALLSVTFW10V20_RF_RCTD 
XI23 VSS VSS TSMC_35 TSMC_36 VDDI VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI33 VSS VSS TSMC_18 TSMC_35 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XXrdtrken TSMC_4 TSMC_1 TSMC_2 TSMC_3 TSMC_5 TSMC_6 TSMC_34 TSMC_19 TSMC_36 
+ TSMC_20 TSMC_21 VDD VDDI VSS S6ALLSVTFW10V20_RF_RDTRKEN 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    16FF_2P_D130_v0d2_x1_for_BL_trk
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk TSMC_1 TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 VDD VSS TSMC_6 TSMC_7 TSMC_8 
MNpg_rp TSMC_3 TSMC_5 TSMC_9 VSS nchpg_8trpsr_mac l=20n nfin=2 m=1 
MNpd_rp TSMC_9 TSMC_1 VSS VSS nchpd_8trpsr_mac l=20n nfin=2 m=1 
MNpg_R TSMC_6 TSMC_8 TSMC_10 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MNpd_R TSMC_10 TSMC_11 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpd_L TSMC_11 TSMC_1 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpg_L TSMC_7 VSS TSMC_11 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MPpu_R TSMC_12 TSMC_11 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
MPpu_L TSMC_11 TSMC_1 TSMC_2 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    16FF_2P_D130_v0d2_x1_for_BL_trk_x2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 TSMC_1 TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 
XI1 TSMC_1 TSMC_3 TSMC_4 TSMC_5 TSMC_7 VDD VSS TSMC_10 TSMC_11 TSMC_12 
+ S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk 
XI0 TSMC_1 TSMC_2 TSMC_4 TSMC_6 TSMC_8 VDD VSS TSMC_9 TSMC_11 TSMC_13 
+ S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RBL_TRK_4X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_D130_ARRAY_RBL_TRK_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 VDD VDDAI 
+ VSS TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 
XI4 VDDAI TSMC_22 TSMC_5 TSMC_6 TSMC_8 TSMC_9 TSMC_12 TSMC_13 VDD VSS 
+ TSMC_23 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
+ S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
XI5 VDDAI TSMC_4 TSMC_22 TSMC_6 TSMC_10 TSMC_11 VSS VSS VDD VSS TSMC_15 
+ TSMC_23 TSMC_17 TSMC_20 TSMC_21 
+ S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WL_TRACK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_WL_TRACK TSMC_1 VSS TSMC_2 TSMC_3 
MMRWL VSS TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MMWWL1 VSS TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MMWWL0q VSS TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RWL_TRK_X2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 VDD VDDAI VSS TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
XI4 TSMC_5 VSS TSMC_5 TSMC_12 S6ALLSVTFW10V20_RF_WL_TRACK 
XI5 TSMC_5 VSS TSMC_5 TSMC_12 S6ALLSVTFW10V20_RF_WL_TRACK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PIN_GCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_PIN_GCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 VSS TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 
XD40 VSS TSMC_77 ndio_mac nfin=2 l=200.0n m=1 
XD39 VSS TSMC_49 ndio_mac nfin=2 l=200.0n m=1 
XD34 VSS TSMC_88 ndio_mac nfin=2 l=200.0n m=1 
XD41 VSS TSMC_78 ndio_mac nfin=2 l=200.0n m=1 
XD5<10> VSS TSMC_12 ndio_mac nfin=2 l=200.0n m=1 
XD5<9> VSS TSMC_13 ndio_mac nfin=2 l=200.0n m=1 
XD5<8> VSS TSMC_14 ndio_mac nfin=2 l=200.0n m=1 
XD5<7> VSS TSMC_15 ndio_mac nfin=2 l=200.0n m=1 
XD5<6> VSS TSMC_16 ndio_mac nfin=2 l=200.0n m=1 
XD5<5> VSS TSMC_17 ndio_mac nfin=2 l=200.0n m=1 
XD5<4> VSS TSMC_18 ndio_mac nfin=2 l=200.0n m=1 
XD5<3> VSS TSMC_19 ndio_mac nfin=2 l=200.0n m=1 
XD5<2> VSS TSMC_20 ndio_mac nfin=2 l=200.0n m=1 
XD5<1> VSS TSMC_21 ndio_mac nfin=2 l=200.0n m=1 
XD5<0> VSS TSMC_22 ndio_mac nfin=2 l=200.0n m=1 
XD8 VSS TSMC_81 ndio_mac nfin=2 l=200.0n m=1 
XD4<10> VSS TSMC_34 ndio_mac nfin=2 l=200.0n m=1 
XD4<9> VSS TSMC_35 ndio_mac nfin=2 l=200.0n m=1 
XD4<8> VSS TSMC_36 ndio_mac nfin=2 l=200.0n m=1 
XD4<7> VSS TSMC_37 ndio_mac nfin=2 l=200.0n m=1 
XD4<6> VSS TSMC_38 ndio_mac nfin=2 l=200.0n m=1 
XD4<5> VSS TSMC_39 ndio_mac nfin=2 l=200.0n m=1 
XD4<4> VSS TSMC_40 ndio_mac nfin=2 l=200.0n m=1 
XD4<3> VSS TSMC_41 ndio_mac nfin=2 l=200.0n m=1 
XD4<2> VSS TSMC_42 ndio_mac nfin=2 l=200.0n m=1 
XD4<1> VSS TSMC_43 ndio_mac nfin=2 l=200.0n m=1 
XD4<0> VSS TSMC_44 ndio_mac nfin=2 l=200.0n m=1 
XD25 VSS TSMC_48 ndio_mac nfin=2 l=200.0n m=1 
XD31<2> VSS TSMC_67 ndio_mac nfin=2 l=200.0n m=1 
XD31<1> VSS TSMC_68 ndio_mac nfin=2 l=200.0n m=1 
XD31<0> VSS TSMC_69 ndio_mac nfin=2 l=200.0n m=1 
XD21 VSS TSMC_92 ndio_mac nfin=2 l=200.0n m=1 
XD35<1> VSS TSMC_51 ndio_mac nfin=2 l=200.0n m=1 
XD35<0> VSS TSMC_52 ndio_mac nfin=2 l=200.0n m=1 
XDdummy<0> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<1> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<2> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<3> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<4> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<5> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD30<2> VSS TSMC_64 ndio_mac nfin=2 l=200.0n m=1 
XD30<1> VSS TSMC_65 ndio_mac nfin=2 l=200.0n m=1 
XD30<0> VSS TSMC_66 ndio_mac nfin=2 l=200.0n m=1 
XD28 VSS TSMC_47 ndio_mac nfin=2 l=200.0n m=1 
XD7 VSS TSMC_76 ndio_mac nfin=2 l=200.0n m=1 
XD2<10> VSS TSMC_23 ndio_mac nfin=2 l=200.0n m=1 
XD2<9> VSS TSMC_24 ndio_mac nfin=2 l=200.0n m=1 
XD2<8> VSS TSMC_25 ndio_mac nfin=2 l=200.0n m=1 
XD2<7> VSS TSMC_26 ndio_mac nfin=2 l=200.0n m=1 
XD2<6> VSS TSMC_27 ndio_mac nfin=2 l=200.0n m=1 
XD2<5> VSS TSMC_28 ndio_mac nfin=2 l=200.0n m=1 
XD2<4> VSS TSMC_29 ndio_mac nfin=2 l=200.0n m=1 
XD2<3> VSS TSMC_30 ndio_mac nfin=2 l=200.0n m=1 
XD2<2> VSS TSMC_31 ndio_mac nfin=2 l=200.0n m=1 
XD2<1> VSS TSMC_32 ndio_mac nfin=2 l=200.0n m=1 
XD2<0> VSS TSMC_33 ndio_mac nfin=2 l=200.0n m=1 
XD3<10> VSS TSMC_1 ndio_mac nfin=2 l=200.0n m=1 
XD3<9> VSS TSMC_2 ndio_mac nfin=2 l=200.0n m=1 
XD3<8> VSS TSMC_3 ndio_mac nfin=2 l=200.0n m=1 
XD3<7> VSS TSMC_4 ndio_mac nfin=2 l=200.0n m=1 
XD3<6> VSS TSMC_5 ndio_mac nfin=2 l=200.0n m=1 
XD3<5> VSS TSMC_6 ndio_mac nfin=2 l=200.0n m=1 
XD3<4> VSS TSMC_7 ndio_mac nfin=2 l=200.0n m=1 
XD3<3> VSS TSMC_8 ndio_mac nfin=2 l=200.0n m=1 
XD3<2> VSS TSMC_9 ndio_mac nfin=2 l=200.0n m=1 
XD3<1> VSS TSMC_10 ndio_mac nfin=2 l=200.0n m=1 
XD3<0> VSS TSMC_11 ndio_mac nfin=2 l=200.0n m=1 
XD0<1> VSS TSMC_71 ndio_mac nfin=2 l=200.0n m=1 
XD0<0> VSS TSMC_72 ndio_mac nfin=2 l=200.0n m=1 
XD24 VSS TSMC_46 ndio_mac nfin=2 l=200.0n m=1 
XD26 VSS TSMC_45 ndio_mac nfin=2 l=200.0n m=1 
XD6 VSS TSMC_50 ndio_mac nfin=2 l=200.0n m=1 
XD9 VSS TSMC_73 ndio_mac nfin=2 l=200.0n m=1 
XD20 VSS TSMC_91 ndio_mac nfin=2 l=200.0n m=1 
XD19 VSS TSMC_74 ndio_mac nfin=2 l=200.0n m=1 
XD38<8> VSS TSMC_53 ndio_mac nfin=2 l=200.0n m=1 
XD38<7> VSS TSMC_54 ndio_mac nfin=2 l=200.0n m=1 
XD38<6> VSS TSMC_55 ndio_mac nfin=2 l=200.0n m=1 
XD38<5> VSS TSMC_56 ndio_mac nfin=2 l=200.0n m=1 
XD38<4> VSS TSMC_57 ndio_mac nfin=2 l=200.0n m=1 
XD38<3> VSS TSMC_58 ndio_mac nfin=2 l=200.0n m=1 
XD38<2> VSS TSMC_59 ndio_mac nfin=2 l=200.0n m=1 
XD38<1> VSS TSMC_60 ndio_mac nfin=2 l=200.0n m=1 
XD38<0> VSS TSMC_61 ndio_mac nfin=2 l=200.0n m=1 
XD37 VSS TSMC_75 ndio_mac nfin=2 l=200.0n m=1 
XD42<1> VSS TSMC_79 ndio_mac nfin=2 l=200.0n m=1 
XD42<0> VSS TSMC_80 ndio_mac nfin=2 l=200.0n m=1 
XD1<1> VSS TSMC_89 ndio_mac nfin=2 l=200.0n m=1 
XD1<0> VSS TSMC_90 ndio_mac nfin=2 l=200.0n m=1 
XD29 VSS TSMC_87 ndio_mac nfin=2 l=200.0n m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    N16_2PRF_BITCELL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_N16_2PRF_BITCELL TSMC_1 TSMC_2 TSMC_3 VDD VSS TSMC_4 
+ TSMC_5 TSMC_6 
MNpg_rp TSMC_2 TSMC_3 TSMC_7 VSS nchpg_8trpsr_mac l=20n nfin=2 m=1 
MNpd_rp TSMC_7 TSMC_8 VSS VSS nchpd_8trpsr_mac l=20n nfin=2 m=1 
MNpd_L TSMC_9 TSMC_8 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpd_R TSMC_8 TSMC_9 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpg_R TSMC_5 TSMC_6 TSMC_8 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MNpg_L TSMC_4 TSMC_6 TSMC_9 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MPpu_L TSMC_9 TSMC_8 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
MPpu_R TSMC_8 TSMC_9 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_4X2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_D130_ARRAY_4X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 VDD VDDAI VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ TSMC_14 TSMC_15 TSMC_16 
XI7 VDDAI TSMC_3 TSMC_7 VDD VSS TSMC_9 TSMC_11 TSMC_15 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
XI6 VDDAI TSMC_4 TSMC_8 VDD VSS TSMC_10 TSMC_12 TSMC_16 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
XI5 VDDAI TSMC_3 TSMC_8 VDD VSS TSMC_9 TSMC_11 TSMC_16 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
XI4 VDDAI TSMC_4 TSMC_7 VDD VSS TSMC_10 TSMC_12 TSMC_15 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
XI3 VDDAI TSMC_4 TSMC_6 VDD VSS TSMC_10 TSMC_12 TSMC_14 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
XI2 VDDAI TSMC_3 TSMC_6 VDD VSS TSMC_9 TSMC_11 TSMC_14 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
XI1 VDDAI TSMC_4 TSMC_5 VDD VSS TSMC_10 TSMC_12 TSMC_13 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
XI0 VDDAI TSMC_3 TSMC_5 VDD VSS TSMC_9 TSMC_11 TSMC_13 
+ S6ALLSVTFW10V20_N16_2PRF_BITCELL 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RBL_TRK_OFF_4X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_D130_ARRAY_RBL_TRK_OFF_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDAI VSS TSMC_12 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
XI2 VDDAI TSMC_4 TSMC_20 TSMC_6 TSMC_10 TSMC_11 VSS VSS VDD VSS TSMC_12 
+ TSMC_21 TSMC_15 TSMC_18 TSMC_19 
+ S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
XI4 VDDAI TSMC_20 TSMC_5 TSMC_6 TSMC_8 TSMC_9 VSS VSS VDD VSS TSMC_21 
+ TSMC_13 TSMC_15 TSMC_16 TSMC_17 
+ S6ALLSVTFW10V20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RWL_TRK_X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X1 TSMC_1 TSMC_2 TSMC_3 VDD VDDAI 
+ VSS TSMC_4 TSMC_5 TSMC_6 TSMC_7 
XI2 TSMC_3 VSS TSMC_3 TSMC_7 S6ALLSVTFW10V20_RF_WL_TRACK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    LIO_PWR_TK_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_LIO_PWR_TK_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI 
+ TSMC_5 
MM_TKPKP3 TSMC_6 TSMC_3 TSMC_7 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP2 TSMC_7 TSMC_3 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP4 TSMC_5 TSMC_4 TSMC_6 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP1 TSMC_6 TSMC_2 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKLIO_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TRKLIO_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS 
MM0 TSMC_3 TSMC_4 VSS VSS nch_lvt_mac l=0.020u nfin=7 m=2 
MM5 TSMC_11 TSMC_9 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_1 TSMC_9 TSMC_11 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_9 TSMC_1 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM8 TSMC_12 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_9 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=2 
MM11 VDD TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_9 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=2 
MM7 TSMC_14 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM13 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM14 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_9 TSMC_1 TSMC_14 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI13 TSMC_5 TSMC_6 TSMC_7 TSMC_10 VDD VDDI TSMC_13 
+ S6ALLSVTFW10V20_LIO_PWR_TK_SVT_V1 
XXpwd0 TSMC_5 TSMC_6 TSMC_7 TSMC_10 VDD VDDI TSMC_13 
+ S6ALLSVTFW10V20_LIO_PWR_TK_SVT_V1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKLIOX2_72_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_TRKLIOX2_72_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 VDD VDDAI VDDI VSS TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 
XI35 VSS VSS TSMC_25 TSMC_26 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI31 VSS VSS TSMC_27 TSMC_28 VDD VDD S6ALLSVTFW10V20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XXtrklio TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_9 TSMC_10 TSMC_11 TSMC_26 TSMC_15 
+ TSMC_18 VDD VDDI VSS S6ALLSVTFW10V20_RF_TRKLIO_SVT_V1 
XI32 TSMC_14 TSMC_1 VSS VSS VDD VDD TSMC_27 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI38 TSMC_28 TSMC_16 VSS VSS VDD VDD TSMC_25 
+ S6ALLSVTFW10V20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    LIO_PWR_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_LIO_PWR_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI 
+ TSMC_5 
MM_PKP3 TSMC_5 TSMC_2 TSMC_6 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_PKP2 TSMC_6 TSMC_2 TSMC_7 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_PKP1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LIO_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_LIO_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 VDD VDDI VSS 
MM4 TSMC_1 TSMC_10 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM8 TSMC_11 TSMC_8 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_1 TSMC_7 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_2 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_2 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_13 TSMC_7 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI0 TSMC_4 TSMC_5 TSMC_6 TSMC_9 VDD VDD TSMC_12 
+ S6ALLSVTFW10V20_LIO_PWR_SVT_V1 
MM2 TSMC_3 TSMC_10 VSS VSS nch_lvt_mac l=0.020u nfin=7 m=2 
XI17 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW10V20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LIOX2_72_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_RF_LIOX2_72_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDAI VDDI VSS 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 
XXlio0 TSMC_9 TSMC_11 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_12 
+ VDD VDDI VSS S6ALLSVTFW10V20_RF_LIO_SVT_V1 
XXlio1 TSMC_8 TSMC_10 TSMC_1 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_12 
+ VDD VDDI VSS S6ALLSVTFW10V20_RF_LIO_SVT_V1 
.ENDS

.SUBCKT ndio_mac PLUS MINUS 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_inv_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_ulvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_inv_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_ulvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nand3_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_lvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nor2_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_ulvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nor2_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_lvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nand2_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_ulvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW10V20_nand2_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS





**** End of leaf cells

.SUBCKT S6ALLSVTFW10V20_PIN_ROW TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 VSS TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 
XPINIO0 TSMC_96 TSMC_210 TSMC_32 TSMC_178 TSMC_64 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO1 TSMC_95 TSMC_209 TSMC_31 TSMC_177 TSMC_63 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO2 TSMC_94 TSMC_208 TSMC_30 TSMC_176 TSMC_62 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO3 TSMC_93 TSMC_207 TSMC_29 TSMC_175 TSMC_61 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO4 TSMC_92 TSMC_206 TSMC_28 TSMC_174 TSMC_60 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO5 TSMC_91 TSMC_205 TSMC_27 TSMC_173 TSMC_59 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO6 TSMC_90 TSMC_204 TSMC_26 TSMC_172 TSMC_58 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO7 TSMC_89 TSMC_203 TSMC_25 TSMC_171 TSMC_57 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO8 TSMC_88 TSMC_202 TSMC_24 TSMC_170 TSMC_56 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO9 TSMC_87 TSMC_201 TSMC_23 TSMC_169 TSMC_55 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO10 TSMC_86 TSMC_200 TSMC_22 TSMC_168 TSMC_54 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO11 TSMC_85 TSMC_199 TSMC_21 TSMC_167 TSMC_53 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO12 TSMC_84 TSMC_198 TSMC_20 TSMC_166 TSMC_52 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO13 TSMC_83 TSMC_197 TSMC_19 TSMC_165 TSMC_51 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO14 TSMC_82 TSMC_196 TSMC_18 TSMC_164 TSMC_50 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO15 TSMC_81 TSMC_195 TSMC_17 TSMC_163 TSMC_49 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO16 TSMC_80 TSMC_194 TSMC_16 TSMC_162 TSMC_48 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO17 TSMC_79 TSMC_193 TSMC_15 TSMC_161 TSMC_47 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO18 TSMC_78 TSMC_192 TSMC_14 TSMC_160 TSMC_46 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO19 TSMC_77 TSMC_191 TSMC_13 TSMC_159 TSMC_45 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO20 TSMC_76 TSMC_190 TSMC_12 TSMC_158 TSMC_44 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO21 TSMC_75 TSMC_189 TSMC_11 TSMC_157 TSMC_43 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO22 TSMC_74 TSMC_188 TSMC_10 TSMC_156 TSMC_42 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO23 TSMC_73 TSMC_187 TSMC_9 TSMC_155 TSMC_41 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO24 TSMC_72 TSMC_186 TSMC_8 TSMC_154 TSMC_40 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO25 TSMC_71 TSMC_185 TSMC_7 TSMC_153 TSMC_39 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO26 TSMC_70 TSMC_184 TSMC_6 TSMC_152 TSMC_38 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO27 TSMC_69 TSMC_183 TSMC_5 TSMC_151 TSMC_37 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO28 TSMC_68 TSMC_182 TSMC_4 TSMC_150 TSMC_36 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO29 TSMC_67 TSMC_181 TSMC_3 TSMC_149 TSMC_35 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO30 TSMC_66 TSMC_180 TSMC_2 TSMC_148 TSMC_34 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINIO31 TSMC_65 TSMC_179 TSMC_1 TSMC_147 TSMC_33 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW10V20_RF_PIN_GIO_MUX2 
XPINCTRL TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_97 TSMC_98 TSMC_99 TSMC_100 
+ TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_136 
+ TSMC_235 TSMC_108 TSMC_121 TSMC_243 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 
+ TSMC_144 TSMC_145 TSMC_253 TSMC_254 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_236 TSMC_129 TSMC_130 TSMC_109 
+ TSMC_233 TSMC_146 TSMC_135 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_134 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_133 VSS TSMC_237 
+ TSMC_131 TSMC_132 TSMC_122 TSMC_234 S6ALLSVTFW10V20_RF_PIN_GCTRL 
.ENDS

.SUBCKT S6ALLSVTFW10V20_GCTRL_GIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 VDDI VDDM VSS TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 
+ TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 
+ TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 
+ TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 
+ TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 
+ TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 
+ TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 
+ TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 
+ TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 
+ TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 
+ TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 
+ TSMC_417 TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 
+ TSMC_425 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 
+ TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 
+ TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 
+ TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 
+ TSMC_473 TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 
+ TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 
+ TSMC_489 TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_504 
+ TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 
+ TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 
+ TSMC_521 TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 
+ TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 
+ TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 
+ TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 
+ TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 TSMC_567 TSMC_568 
+ TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 TSMC_578 TSMC_579 TSMC_580 TSMC_581 TSMC_582 TSMC_583 
XGIO_MUX0 TSMC_34 TSMC_66 TSMC_129 TSMC_130 TSMC_550 TSMC_582 TSMC_584 TSMC_178 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_454 TSMC_518 
+ TSMC_486 TSMC_282 TSMC_283 TSMC_346 TSMC_347 TSMC_382 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX1 TSMC_33 TSMC_65 TSMC_127 TSMC_128 TSMC_549 TSMC_581 TSMC_584 TSMC_177 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_453 TSMC_517 
+ TSMC_485 TSMC_280 TSMC_281 TSMC_344 TSMC_345 TSMC_381 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX2 TSMC_32 TSMC_64 TSMC_125 TSMC_126 TSMC_548 TSMC_580 TSMC_584 TSMC_176 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_452 TSMC_516 
+ TSMC_484 TSMC_278 TSMC_279 TSMC_342 TSMC_343 TSMC_380 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX3 TSMC_31 TSMC_63 TSMC_123 TSMC_124 TSMC_547 TSMC_579 TSMC_584 TSMC_175 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_451 TSMC_515 
+ TSMC_483 TSMC_276 TSMC_277 TSMC_340 TSMC_341 TSMC_379 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX4 TSMC_30 TSMC_62 TSMC_121 TSMC_122 TSMC_546 TSMC_578 TSMC_584 TSMC_174 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_450 TSMC_514 
+ TSMC_482 TSMC_274 TSMC_275 TSMC_338 TSMC_339 TSMC_378 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX5 TSMC_29 TSMC_61 TSMC_119 TSMC_120 TSMC_545 TSMC_577 TSMC_584 TSMC_173 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_449 TSMC_513 
+ TSMC_481 TSMC_272 TSMC_273 TSMC_336 TSMC_337 TSMC_377 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX6 TSMC_28 TSMC_60 TSMC_117 TSMC_118 TSMC_544 TSMC_576 TSMC_584 TSMC_172 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_448 TSMC_512 
+ TSMC_480 TSMC_270 TSMC_271 TSMC_334 TSMC_335 TSMC_376 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX7 TSMC_27 TSMC_59 TSMC_115 TSMC_116 TSMC_543 TSMC_575 TSMC_584 TSMC_171 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_447 TSMC_511 
+ TSMC_479 TSMC_268 TSMC_269 TSMC_332 TSMC_333 TSMC_375 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX8 TSMC_26 TSMC_58 TSMC_113 TSMC_114 TSMC_542 TSMC_574 TSMC_584 TSMC_170 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_446 TSMC_510 
+ TSMC_478 TSMC_266 TSMC_267 TSMC_330 TSMC_331 TSMC_374 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX9 TSMC_25 TSMC_57 TSMC_111 TSMC_112 TSMC_541 TSMC_573 TSMC_584 TSMC_169 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_445 TSMC_509 
+ TSMC_477 TSMC_264 TSMC_265 TSMC_328 TSMC_329 TSMC_373 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX10 TSMC_24 TSMC_56 TSMC_109 TSMC_110 TSMC_540 TSMC_572 TSMC_584 
+ TSMC_168 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_444 
+ TSMC_508 TSMC_476 TSMC_262 TSMC_263 TSMC_326 TSMC_327 TSMC_372 
+ TSMC_588 TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 
+ TSMC_592 S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX11 TSMC_23 TSMC_55 TSMC_107 TSMC_108 TSMC_539 TSMC_571 TSMC_584 
+ TSMC_167 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_443 
+ TSMC_507 TSMC_475 TSMC_260 TSMC_261 TSMC_324 TSMC_325 TSMC_371 
+ TSMC_588 TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 
+ TSMC_590 S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX12 TSMC_22 TSMC_54 TSMC_105 TSMC_106 TSMC_538 TSMC_570 TSMC_584 
+ TSMC_166 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_442 
+ TSMC_506 TSMC_474 TSMC_258 TSMC_259 TSMC_322 TSMC_323 TSMC_370 
+ TSMC_588 TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 
+ TSMC_592 S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX13 TSMC_21 TSMC_53 TSMC_103 TSMC_104 TSMC_537 TSMC_569 TSMC_584 
+ TSMC_165 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_441 
+ TSMC_505 TSMC_473 TSMC_256 TSMC_257 TSMC_320 TSMC_321 TSMC_369 
+ TSMC_588 TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 
+ TSMC_590 S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX14 TSMC_20 TSMC_52 TSMC_101 TSMC_102 TSMC_536 TSMC_568 TSMC_584 
+ TSMC_164 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_440 
+ TSMC_504 TSMC_472 TSMC_254 TSMC_255 TSMC_318 TSMC_319 TSMC_368 
+ TSMC_588 TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 
+ TSMC_592 S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX15 TSMC_19 TSMC_51 TSMC_99 TSMC_100 TSMC_535 TSMC_567 TSMC_584 
+ TSMC_163 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_439 TSMC_503 
+ TSMC_471 TSMC_252 TSMC_253 TSMC_316 TSMC_317 TSMC_367 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX16 TSMC_18 TSMC_50 TSMC_97 TSMC_98 TSMC_534 TSMC_566 TSMC_584 
+ TSMC_162 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_438 TSMC_502 
+ TSMC_470 TSMC_250 TSMC_251 TSMC_314 TSMC_315 TSMC_366 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX17 TSMC_17 TSMC_49 TSMC_95 TSMC_96 TSMC_533 TSMC_565 TSMC_584 
+ TSMC_161 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_437 TSMC_501 
+ TSMC_469 TSMC_248 TSMC_249 TSMC_312 TSMC_313 TSMC_365 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX18 TSMC_16 TSMC_48 TSMC_93 TSMC_94 TSMC_532 TSMC_564 TSMC_584 
+ TSMC_160 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_436 TSMC_500 
+ TSMC_468 TSMC_246 TSMC_247 TSMC_310 TSMC_311 TSMC_364 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX19 TSMC_15 TSMC_47 TSMC_91 TSMC_92 TSMC_531 TSMC_563 TSMC_584 
+ TSMC_159 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_435 TSMC_499 
+ TSMC_467 TSMC_244 TSMC_245 TSMC_308 TSMC_309 TSMC_363 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX20 TSMC_14 TSMC_46 TSMC_89 TSMC_90 TSMC_530 TSMC_562 TSMC_584 
+ TSMC_158 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_434 TSMC_498 
+ TSMC_466 TSMC_242 TSMC_243 TSMC_306 TSMC_307 TSMC_362 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX21 TSMC_13 TSMC_45 TSMC_87 TSMC_88 TSMC_529 TSMC_561 TSMC_584 
+ TSMC_157 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_433 TSMC_497 
+ TSMC_465 TSMC_240 TSMC_241 TSMC_304 TSMC_305 TSMC_361 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX22 TSMC_12 TSMC_44 TSMC_85 TSMC_86 TSMC_528 TSMC_560 TSMC_584 
+ TSMC_156 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_432 TSMC_496 
+ TSMC_464 TSMC_238 TSMC_239 TSMC_302 TSMC_303 TSMC_360 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX23 TSMC_11 TSMC_43 TSMC_83 TSMC_84 TSMC_527 TSMC_559 TSMC_584 
+ TSMC_155 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_431 TSMC_495 
+ TSMC_463 TSMC_236 TSMC_237 TSMC_300 TSMC_301 TSMC_359 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX24 TSMC_10 TSMC_42 TSMC_81 TSMC_82 TSMC_526 TSMC_558 TSMC_584 
+ TSMC_154 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_430 TSMC_494 
+ TSMC_462 TSMC_234 TSMC_235 TSMC_298 TSMC_299 TSMC_358 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX25 TSMC_9 TSMC_41 TSMC_79 TSMC_80 TSMC_525 TSMC_557 TSMC_584 
+ TSMC_153 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_429 TSMC_493 
+ TSMC_461 TSMC_232 TSMC_233 TSMC_296 TSMC_297 TSMC_357 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX26 TSMC_8 TSMC_40 TSMC_77 TSMC_78 TSMC_524 TSMC_556 TSMC_584 
+ TSMC_152 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_428 TSMC_492 
+ TSMC_460 TSMC_230 TSMC_231 TSMC_294 TSMC_295 TSMC_356 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX27 TSMC_7 TSMC_39 TSMC_75 TSMC_76 TSMC_523 TSMC_555 TSMC_584 
+ TSMC_151 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_427 TSMC_491 
+ TSMC_459 TSMC_228 TSMC_229 TSMC_292 TSMC_293 TSMC_355 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX28 TSMC_6 TSMC_38 TSMC_73 TSMC_74 TSMC_522 TSMC_554 TSMC_584 
+ TSMC_150 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_426 TSMC_490 
+ TSMC_458 TSMC_226 TSMC_227 TSMC_290 TSMC_291 TSMC_354 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX29 TSMC_5 TSMC_37 TSMC_71 TSMC_72 TSMC_521 TSMC_553 TSMC_584 
+ TSMC_149 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_425 TSMC_489 
+ TSMC_457 TSMC_224 TSMC_225 TSMC_288 TSMC_289 TSMC_353 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX30 TSMC_4 TSMC_36 TSMC_69 TSMC_70 TSMC_520 TSMC_552 TSMC_584 
+ TSMC_148 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_424 TSMC_488 
+ TSMC_456 TSMC_222 TSMC_223 TSMC_286 TSMC_287 TSMC_352 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_GIOM2 
XGIO_MUX31 TSMC_3 TSMC_35 TSMC_67 TSMC_68 TSMC_519 TSMC_551 TSMC_584 
+ TSMC_147 TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_423 TSMC_487 
+ TSMC_455 TSMC_220 TSMC_221 TSMC_284 TSMC_285 TSMC_351 TSMC_588 
+ TSMC_418 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_589 TSMC_590 
+ S6ALLSVTFW10V20_RF_GIOM2 
XTRKGIOL TSMC_584 TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_216 VDDM VDDI VSS TSMC_599 TSMC_600 
+ TSMC_144 TSMC_348 TSMC_349 TSMC_145 TSMC_588 TSMC_418 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_589 TSMC_590 TSMC_591 
+ TSMC_592 S6ALLSVTFW10V20_RF_TRKGIOWR 
XTRKGIOR TSMC_606 TSMC_607 TSMC_608 TSMC_131 TSMC_217 TSMC_217 TSMC_584 
+ TSMC_179 TSMC_180 TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 
+ TSMC_598 TSMC_585 TSMC_586 TSMC_587 TSMC_609 TSMC_217 TSMC_216 VDDM 
+ VDDI VSS TSMC_415 TSMC_610 TSMC_588 TSMC_418 TSMC_602 TSMC_603 
+ TSMC_604 TSMC_605 TSMC_589 TSMC_590 TSMC_591 TSMC_592 
+ S6ALLSVTFW10V20_RF_TRKGIORD 
XGCTRL TSMC_1 TSMC_2 TSMC_420 TSMC_611 TSMC_421 TSMC_422 TSMC_419 TSMC_132 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_216 TSMC_216 TSMC_612 
+ TSMC_217 TSMC_217 TSMC_613 TSMC_614 TSMC_416 TSMC_146 TSMC_584 TSMC_417 
+ TSMC_615 TSMC_616 TSMC_615 TSMC_616 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_617 TSMC_618 TSMC_612 TSMC_619 
+ TSMC_620 TSMC_613 TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 
+ TSMC_598 TSMC_585 TSMC_586 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 
+ TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_587 TSMC_203 TSMC_609 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_583 TSMC_217 TSMC_216 
+ TSMC_218 TSMC_219 VDDM VDDI VSS TSMC_350 TSMC_383 TSMC_384 TSMC_385 
+ TSMC_588 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 
+ TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 
+ TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_418 TSMC_601 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_602 TSMC_603 TSMC_604 TSMC_605 
+ TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_621 TSMC_622 TSMC_615 
+ TSMC_616 S6ALLSVTFW10V20_RF_GCTRL 
.ENDS

.SUBCKT S6ALLSVTFW10V20_ROW_TRACKING TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 VDDM 
+ VDDAI VDDI VSS TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 
XTRKROW0 TSMC_191 TSMC_192 TSMC_200 TSMC_201 TSMC_197 VDDM VDDAI VSS TSMC_63 
+ TSMC_64 TSMC_127 TSMC_128 TSMC_202 TSMC_203 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW1 TSMC_189 TSMC_190 TSMC_204 TSMC_205 TSMC_197 VDDM VDDAI VSS TSMC_61 
+ TSMC_62 TSMC_125 TSMC_126 TSMC_206 TSMC_207 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW2 TSMC_187 TSMC_188 TSMC_208 TSMC_209 TSMC_197 VDDM VDDAI VSS TSMC_59 
+ TSMC_60 TSMC_123 TSMC_124 TSMC_210 TSMC_211 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW3 TSMC_185 TSMC_186 TSMC_212 TSMC_213 TSMC_197 VDDM VDDAI VSS TSMC_57 
+ TSMC_58 TSMC_121 TSMC_122 TSMC_214 TSMC_215 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW4 TSMC_183 TSMC_184 TSMC_216 TSMC_217 TSMC_197 VDDM VDDAI VSS TSMC_55 
+ TSMC_56 TSMC_119 TSMC_120 TSMC_218 TSMC_219 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW5 TSMC_181 TSMC_182 TSMC_220 TSMC_221 TSMC_197 VDDM VDDAI VSS TSMC_53 
+ TSMC_54 TSMC_117 TSMC_118 TSMC_222 TSMC_223 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW6 TSMC_179 TSMC_180 TSMC_224 TSMC_225 TSMC_197 VDDM VDDAI VSS TSMC_51 
+ TSMC_52 TSMC_115 TSMC_116 TSMC_226 TSMC_227 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW7 TSMC_177 TSMC_178 TSMC_228 TSMC_229 TSMC_197 VDDM VDDAI VSS TSMC_49 
+ TSMC_50 TSMC_113 TSMC_114 TSMC_230 TSMC_231 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW8 TSMC_175 TSMC_176 TSMC_232 TSMC_233 TSMC_197 VDDM VDDAI VSS TSMC_47 
+ TSMC_48 TSMC_111 TSMC_112 TSMC_234 TSMC_235 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW9 TSMC_173 TSMC_174 TSMC_236 TSMC_237 TSMC_197 VDDM VDDAI VSS TSMC_45 
+ TSMC_46 TSMC_109 TSMC_110 TSMC_238 TSMC_239 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW10 TSMC_171 TSMC_172 TSMC_240 TSMC_241 TSMC_197 VDDM VDDAI VSS TSMC_43 
+ TSMC_44 TSMC_107 TSMC_108 TSMC_242 TSMC_243 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW11 TSMC_169 TSMC_170 TSMC_244 TSMC_245 TSMC_197 VDDM VDDAI VSS TSMC_41 
+ TSMC_42 TSMC_105 TSMC_106 TSMC_246 TSMC_247 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW12 TSMC_167 TSMC_168 TSMC_248 TSMC_249 TSMC_197 VDDM VDDAI VSS TSMC_39 
+ TSMC_40 TSMC_103 TSMC_104 TSMC_250 TSMC_251 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW13 TSMC_165 TSMC_166 TSMC_252 TSMC_253 TSMC_197 VDDM VDDAI VSS TSMC_37 
+ TSMC_38 TSMC_101 TSMC_102 TSMC_254 TSMC_255 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW14 TSMC_163 TSMC_164 TSMC_256 TSMC_257 TSMC_197 VDDM VDDAI VSS TSMC_35 
+ TSMC_36 TSMC_99 TSMC_100 TSMC_258 TSMC_259 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW15 TSMC_161 TSMC_162 TSMC_260 TSMC_261 TSMC_197 VDDM VDDAI VSS TSMC_33 
+ TSMC_34 TSMC_97 TSMC_98 TSMC_262 TSMC_263 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW16 TSMC_159 TSMC_160 TSMC_264 TSMC_265 TSMC_197 VDDM VDDAI VSS TSMC_31 
+ TSMC_32 TSMC_95 TSMC_96 TSMC_266 TSMC_267 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW17 TSMC_157 TSMC_158 TSMC_268 TSMC_269 TSMC_197 VDDM VDDAI VSS TSMC_29 
+ TSMC_30 TSMC_93 TSMC_94 TSMC_270 TSMC_271 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW18 TSMC_155 TSMC_156 TSMC_272 TSMC_273 TSMC_197 VDDM VDDAI VSS TSMC_27 
+ TSMC_28 TSMC_91 TSMC_92 TSMC_274 TSMC_275 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW19 TSMC_153 TSMC_154 TSMC_276 TSMC_277 TSMC_197 VDDM VDDAI VSS TSMC_25 
+ TSMC_26 TSMC_89 TSMC_90 TSMC_278 TSMC_279 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW20 TSMC_151 TSMC_152 TSMC_280 TSMC_281 TSMC_197 VDDM VDDAI VSS TSMC_23 
+ TSMC_24 TSMC_87 TSMC_88 TSMC_282 TSMC_283 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW21 TSMC_149 TSMC_150 TSMC_284 TSMC_285 TSMC_197 VDDM VDDAI VSS TSMC_21 
+ TSMC_22 TSMC_85 TSMC_86 TSMC_286 TSMC_287 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW22 TSMC_147 TSMC_148 TSMC_288 TSMC_289 TSMC_197 VDDM VDDAI VSS TSMC_19 
+ TSMC_20 TSMC_83 TSMC_84 TSMC_290 TSMC_291 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW23 TSMC_145 TSMC_146 TSMC_292 TSMC_293 TSMC_197 VDDM VDDAI VSS TSMC_17 
+ TSMC_18 TSMC_81 TSMC_82 TSMC_294 TSMC_295 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW24 TSMC_143 TSMC_144 TSMC_296 TSMC_297 TSMC_197 VDDM VDDAI VSS TSMC_15 
+ TSMC_16 TSMC_79 TSMC_80 TSMC_298 TSMC_299 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW25 TSMC_141 TSMC_142 TSMC_300 TSMC_301 TSMC_197 VDDM VDDAI VSS TSMC_13 
+ TSMC_14 TSMC_77 TSMC_78 TSMC_302 TSMC_303 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW26 TSMC_139 TSMC_140 TSMC_304 TSMC_305 TSMC_197 VDDM VDDAI VSS TSMC_11 
+ TSMC_12 TSMC_75 TSMC_76 TSMC_306 TSMC_307 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW27 TSMC_137 TSMC_138 TSMC_308 TSMC_309 TSMC_197 VDDM VDDAI VSS TSMC_9 
+ TSMC_10 TSMC_73 TSMC_74 TSMC_310 TSMC_311 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW28 TSMC_135 TSMC_136 TSMC_312 TSMC_313 TSMC_197 VDDM VDDAI VSS TSMC_7 
+ TSMC_8 TSMC_71 TSMC_72 TSMC_314 TSMC_315 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW29 TSMC_133 TSMC_134 TSMC_316 TSMC_317 TSMC_197 VDDM VDDAI VSS TSMC_5 
+ TSMC_6 TSMC_69 TSMC_70 TSMC_318 TSMC_319 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW30 TSMC_131 TSMC_132 TSMC_320 TSMC_321 TSMC_197 VDDM VDDAI VSS TSMC_3 
+ TSMC_4 TSMC_67 TSMC_68 TSMC_322 TSMC_323 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROW31 TSMC_129 TSMC_130 TSMC_324 TSMC_325 TSMC_197 VDDM VDDAI VSS TSMC_1 
+ TSMC_2 TSMC_65 TSMC_66 TSMC_326 TSMC_327 VSS 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XTRKROWL TSMC_328 TSMC_329 TSMC_197 VDDM VDDAI VSS TSMC_198 TSMC_330 
+ TSMC_331 VSS S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X1 
XTRKROWR TSMC_193 TSMC_332 TSMC_197 VDDM VDDAI VSS TSMC_199 TSMC_333 
+ TSMC_334 VSS S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X1 
XTRKCTRL TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 
+ TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_196 TSMC_194 TSMC_195 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 
+ TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 
+ TSMC_360 TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_197 VDDM VDDI VSS TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 
+ TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_377 TSMC_378 TSMC_379 
+ TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 
+ S6ALLSVTFW10V20_RF_TRKCTRL 
.ENDS

.SUBCKT S6ALLSVTFW10V20_ARY4ROW TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 VDDM VDDAI 
+ VDDI VSS TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 
+ TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 
+ TSMC_296 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
XCOL0 TSMC_63 TSMC_64 TSMC_127 TSMC_128 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_191 TSMC_192 TSMC_255 TSMC_256 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL1 TSMC_61 TSMC_62 TSMC_125 TSMC_126 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_189 TSMC_190 TSMC_253 TSMC_254 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL2 TSMC_59 TSMC_60 TSMC_123 TSMC_124 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_187 TSMC_188 TSMC_251 TSMC_252 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL3 TSMC_57 TSMC_58 TSMC_121 TSMC_122 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_185 TSMC_186 TSMC_249 TSMC_250 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL4 TSMC_55 TSMC_56 TSMC_119 TSMC_120 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_183 TSMC_184 TSMC_247 TSMC_248 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL5 TSMC_53 TSMC_54 TSMC_117 TSMC_118 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_181 TSMC_182 TSMC_245 TSMC_246 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL6 TSMC_51 TSMC_52 TSMC_115 TSMC_116 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_179 TSMC_180 TSMC_243 TSMC_244 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL7 TSMC_49 TSMC_50 TSMC_113 TSMC_114 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_177 TSMC_178 TSMC_241 TSMC_242 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL8 TSMC_47 TSMC_48 TSMC_111 TSMC_112 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_175 TSMC_176 TSMC_239 TSMC_240 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL9 TSMC_45 TSMC_46 TSMC_109 TSMC_110 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_173 TSMC_174 TSMC_237 TSMC_238 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL10 TSMC_43 TSMC_44 TSMC_107 TSMC_108 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_171 TSMC_172 TSMC_235 TSMC_236 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL11 TSMC_41 TSMC_42 TSMC_105 TSMC_106 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_169 TSMC_170 TSMC_233 TSMC_234 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL12 TSMC_39 TSMC_40 TSMC_103 TSMC_104 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_167 TSMC_168 TSMC_231 TSMC_232 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL13 TSMC_37 TSMC_38 TSMC_101 TSMC_102 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_165 TSMC_166 TSMC_229 TSMC_230 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL14 TSMC_35 TSMC_36 TSMC_99 TSMC_100 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ VDDM VDDAI VSS TSMC_163 TSMC_164 TSMC_227 TSMC_228 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL15 TSMC_33 TSMC_34 TSMC_97 TSMC_98 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_161 TSMC_162 TSMC_225 TSMC_226 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL16 TSMC_31 TSMC_32 TSMC_95 TSMC_96 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_159 TSMC_160 TSMC_223 TSMC_224 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL17 TSMC_29 TSMC_30 TSMC_93 TSMC_94 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_157 TSMC_158 TSMC_221 TSMC_222 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL18 TSMC_27 TSMC_28 TSMC_91 TSMC_92 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_155 TSMC_156 TSMC_219 TSMC_220 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL19 TSMC_25 TSMC_26 TSMC_89 TSMC_90 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_153 TSMC_154 TSMC_217 TSMC_218 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL20 TSMC_23 TSMC_24 TSMC_87 TSMC_88 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_151 TSMC_152 TSMC_215 TSMC_216 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL21 TSMC_21 TSMC_22 TSMC_85 TSMC_86 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_149 TSMC_150 TSMC_213 TSMC_214 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL22 TSMC_19 TSMC_20 TSMC_83 TSMC_84 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_147 TSMC_148 TSMC_211 TSMC_212 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL23 TSMC_17 TSMC_18 TSMC_81 TSMC_82 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_145 TSMC_146 TSMC_209 TSMC_210 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL24 TSMC_15 TSMC_16 TSMC_79 TSMC_80 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_143 TSMC_144 TSMC_207 TSMC_208 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL25 TSMC_13 TSMC_14 TSMC_77 TSMC_78 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_141 TSMC_142 TSMC_205 TSMC_206 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL26 TSMC_11 TSMC_12 TSMC_75 TSMC_76 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_139 TSMC_140 TSMC_203 TSMC_204 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL27 TSMC_9 TSMC_10 TSMC_73 TSMC_74 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_137 TSMC_138 TSMC_201 TSMC_202 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL28 TSMC_7 TSMC_8 TSMC_71 TSMC_72 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_135 TSMC_136 TSMC_199 TSMC_200 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL29 TSMC_5 TSMC_6 TSMC_69 TSMC_70 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_133 TSMC_134 TSMC_197 TSMC_198 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL30 TSMC_3 TSMC_4 TSMC_67 TSMC_68 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_131 TSMC_132 TSMC_195 TSMC_196 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL31 TSMC_1 TSMC_2 TSMC_65 TSMC_66 TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM 
+ VDDAI VSS TSMC_129 TSMC_130 TSMC_193 TSMC_194 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XTRKL TSMC_257 TSMC_320 TSMC_321 TSMC_308 TSMC_309 TSMC_258 TSMC_258 
+ TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM VDDAI VSS TSMC_304 TSMC_305 VSS 
+ TSMC_259 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ S6ALLSVTFW10V20_D130_ARRAY_RBL_TRK_OFF_4X1 
XTRKR TSMC_260 TSMC_322 TSMC_323 TSMC_310 TSMC_311 TSMC_258 TSMC_258 
+ TSMC_312 TSMC_313 TSMC_314 TSMC_315 VDDM VDDAI VSS TSMC_306 TSMC_307 VSS 
+ TSMC_261 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ S6ALLSVTFW10V20_D130_ARRAY_RBL_TRK_OFF_4X1 
XDEC TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 
+ TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 
+ TSMC_339 TSMC_340 TSMC_262 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_280 VDDM VDDI VDDI VSS TSMC_281 
+ TSMC_282 TSMC_283 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 
+ TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 
+ TSMC_295 TSMC_296 TSMC_297 TSMC_298 TSMC_299 TSMC_316 TSMC_317 TSMC_318 
+ TSMC_319 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ S6ALLSVTFW10V20_RF_XDEC4 
.ENDS

.SUBCKT S6ALLSVTFW10V20_ARY4ROW_TK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 VDDM VDDAI 
+ VDDI VSS TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 
+ TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 
+ TSMC_296 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
+ TSMC_312 TSMC_313 
XCOL0 TSMC_63 TSMC_64 TSMC_127 TSMC_128 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_191 TSMC_192 TSMC_255 TSMC_256 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL1 TSMC_61 TSMC_62 TSMC_125 TSMC_126 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_189 TSMC_190 TSMC_253 TSMC_254 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL2 TSMC_59 TSMC_60 TSMC_123 TSMC_124 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_187 TSMC_188 TSMC_251 TSMC_252 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL3 TSMC_57 TSMC_58 TSMC_121 TSMC_122 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_185 TSMC_186 TSMC_249 TSMC_250 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL4 TSMC_55 TSMC_56 TSMC_119 TSMC_120 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_183 TSMC_184 TSMC_247 TSMC_248 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL5 TSMC_53 TSMC_54 TSMC_117 TSMC_118 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_181 TSMC_182 TSMC_245 TSMC_246 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL6 TSMC_51 TSMC_52 TSMC_115 TSMC_116 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_179 TSMC_180 TSMC_243 TSMC_244 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL7 TSMC_49 TSMC_50 TSMC_113 TSMC_114 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_177 TSMC_178 TSMC_241 TSMC_242 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL8 TSMC_47 TSMC_48 TSMC_111 TSMC_112 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_175 TSMC_176 TSMC_239 TSMC_240 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL9 TSMC_45 TSMC_46 TSMC_109 TSMC_110 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_173 TSMC_174 TSMC_237 TSMC_238 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL10 TSMC_43 TSMC_44 TSMC_107 TSMC_108 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_171 TSMC_172 TSMC_235 TSMC_236 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL11 TSMC_41 TSMC_42 TSMC_105 TSMC_106 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_169 TSMC_170 TSMC_233 TSMC_234 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL12 TSMC_39 TSMC_40 TSMC_103 TSMC_104 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_167 TSMC_168 TSMC_231 TSMC_232 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL13 TSMC_37 TSMC_38 TSMC_101 TSMC_102 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_165 TSMC_166 TSMC_229 TSMC_230 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL14 TSMC_35 TSMC_36 TSMC_99 TSMC_100 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ VDDM VDDAI VSS TSMC_163 TSMC_164 TSMC_227 TSMC_228 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL15 TSMC_33 TSMC_34 TSMC_97 TSMC_98 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_161 TSMC_162 TSMC_225 TSMC_226 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL16 TSMC_31 TSMC_32 TSMC_95 TSMC_96 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_159 TSMC_160 TSMC_223 TSMC_224 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL17 TSMC_29 TSMC_30 TSMC_93 TSMC_94 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_157 TSMC_158 TSMC_221 TSMC_222 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL18 TSMC_27 TSMC_28 TSMC_91 TSMC_92 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_155 TSMC_156 TSMC_219 TSMC_220 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL19 TSMC_25 TSMC_26 TSMC_89 TSMC_90 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_153 TSMC_154 TSMC_217 TSMC_218 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL20 TSMC_23 TSMC_24 TSMC_87 TSMC_88 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_151 TSMC_152 TSMC_215 TSMC_216 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL21 TSMC_21 TSMC_22 TSMC_85 TSMC_86 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_149 TSMC_150 TSMC_213 TSMC_214 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL22 TSMC_19 TSMC_20 TSMC_83 TSMC_84 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_147 TSMC_148 TSMC_211 TSMC_212 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL23 TSMC_17 TSMC_18 TSMC_81 TSMC_82 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_145 TSMC_146 TSMC_209 TSMC_210 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL24 TSMC_15 TSMC_16 TSMC_79 TSMC_80 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_143 TSMC_144 TSMC_207 TSMC_208 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL25 TSMC_13 TSMC_14 TSMC_77 TSMC_78 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_141 TSMC_142 TSMC_205 TSMC_206 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL26 TSMC_11 TSMC_12 TSMC_75 TSMC_76 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_139 TSMC_140 TSMC_203 TSMC_204 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL27 TSMC_9 TSMC_10 TSMC_73 TSMC_74 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_137 TSMC_138 TSMC_201 TSMC_202 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL28 TSMC_7 TSMC_8 TSMC_71 TSMC_72 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_135 TSMC_136 TSMC_199 TSMC_200 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL29 TSMC_5 TSMC_6 TSMC_69 TSMC_70 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_133 TSMC_134 TSMC_197 TSMC_198 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL30 TSMC_3 TSMC_4 TSMC_67 TSMC_68 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_131 TSMC_132 TSMC_195 TSMC_196 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XCOL31 TSMC_1 TSMC_2 TSMC_65 TSMC_66 TSMC_314 TSMC_315 TSMC_316 TSMC_317 VDDM 
+ VDDAI VSS TSMC_129 TSMC_130 TSMC_193 TSMC_194 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_4X2 
XTRKL TSMC_257 TSMC_322 TSMC_323 TSMC_310 TSMC_311 TSMC_258 TSMC_258 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_308 TSMC_308 VDDM VDDAI VSS VSS 
+ TSMC_304 TSMC_305 TSMC_259 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_RBL_TRK_4X1 
XTRKR TSMC_324 TSMC_325 TSMC_326 TSMC_312 TSMC_313 TSMC_258 TSMC_258 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_309 TSMC_309 VDDM VDDAI VSS VSS 
+ TSMC_306 TSMC_307 TSMC_261 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 S6ALLSVTFW10V20_D130_ARRAY_RBL_TRK_4X1 
XDEC TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 
+ TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 
+ TSMC_342 TSMC_343 TSMC_262 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_314 
+ TSMC_315 TSMC_316 TSMC_317 TSMC_280 VDDM VDDI VDDI VSS TSMC_281 
+ TSMC_282 TSMC_283 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 
+ TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 
+ TSMC_295 TSMC_296 TSMC_297 TSMC_298 TSMC_299 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ S6ALLSVTFW10V20_RF_XDEC4 
.ENDS

.SUBCKT S6ALLSVTFW10V20_LIO_LCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 
+ TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 
+ TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 VDDM VDDI VDDAI VSS 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 
+ TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 
+ TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 
+ TSMC_400 TSMC_401 
XLIO0 TSMC_63 TSMC_64 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_127 
+ TSMC_128 TSMC_191 TSMC_192 TSMC_373 VDDM VDDAI VDDI VSS TSMC_255 
+ TSMC_256 TSMC_319 TSMC_320 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO1 TSMC_61 TSMC_62 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_125 
+ TSMC_126 TSMC_189 TSMC_190 TSMC_373 VDDM VDDAI VDDI VSS TSMC_253 
+ TSMC_254 TSMC_317 TSMC_318 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO2 TSMC_59 TSMC_60 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_123 
+ TSMC_124 TSMC_187 TSMC_188 TSMC_373 VDDM VDDAI VDDI VSS TSMC_251 
+ TSMC_252 TSMC_315 TSMC_316 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO3 TSMC_57 TSMC_58 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_121 
+ TSMC_122 TSMC_185 TSMC_186 TSMC_373 VDDM VDDAI VDDI VSS TSMC_249 
+ TSMC_250 TSMC_313 TSMC_314 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO4 TSMC_55 TSMC_56 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_119 
+ TSMC_120 TSMC_183 TSMC_184 TSMC_373 VDDM VDDAI VDDI VSS TSMC_247 
+ TSMC_248 TSMC_311 TSMC_312 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO5 TSMC_53 TSMC_54 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_117 
+ TSMC_118 TSMC_181 TSMC_182 TSMC_373 VDDM VDDAI VDDI VSS TSMC_245 
+ TSMC_246 TSMC_309 TSMC_310 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO6 TSMC_51 TSMC_52 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_115 
+ TSMC_116 TSMC_179 TSMC_180 TSMC_373 VDDM VDDAI VDDI VSS TSMC_243 
+ TSMC_244 TSMC_307 TSMC_308 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO7 TSMC_49 TSMC_50 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_113 
+ TSMC_114 TSMC_177 TSMC_178 TSMC_373 VDDM VDDAI VDDI VSS TSMC_241 
+ TSMC_242 TSMC_305 TSMC_306 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO8 TSMC_47 TSMC_48 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_111 
+ TSMC_112 TSMC_175 TSMC_176 TSMC_373 VDDM VDDAI VDDI VSS TSMC_239 
+ TSMC_240 TSMC_303 TSMC_304 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO9 TSMC_45 TSMC_46 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_109 
+ TSMC_110 TSMC_173 TSMC_174 TSMC_373 VDDM VDDAI VDDI VSS TSMC_237 
+ TSMC_238 TSMC_301 TSMC_302 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO10 TSMC_43 TSMC_44 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_107 TSMC_108 TSMC_171 TSMC_172 TSMC_373 VDDM VDDAI VDDI VSS TSMC_235 
+ TSMC_236 TSMC_299 TSMC_300 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO11 TSMC_41 TSMC_42 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_105 TSMC_106 TSMC_169 TSMC_170 TSMC_373 VDDM VDDAI VDDI VSS TSMC_233 
+ TSMC_234 TSMC_297 TSMC_298 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO12 TSMC_39 TSMC_40 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_103 TSMC_104 TSMC_167 TSMC_168 TSMC_373 VDDM VDDAI VDDI VSS TSMC_231 
+ TSMC_232 TSMC_295 TSMC_296 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO13 TSMC_37 TSMC_38 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_101 TSMC_102 TSMC_165 TSMC_166 TSMC_373 VDDM VDDAI VDDI VSS TSMC_229 
+ TSMC_230 TSMC_293 TSMC_294 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO14 TSMC_35 TSMC_36 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_99 TSMC_100 TSMC_163 TSMC_164 TSMC_373 VDDM VDDAI VDDI VSS TSMC_227 
+ TSMC_228 TSMC_291 TSMC_292 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO15 TSMC_33 TSMC_34 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_97 TSMC_98 TSMC_161 TSMC_162 TSMC_373 VDDM VDDAI VDDI VSS TSMC_225 
+ TSMC_226 TSMC_289 TSMC_290 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO16 TSMC_31 TSMC_32 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_95 TSMC_96 TSMC_159 TSMC_160 TSMC_373 VDDM VDDAI VDDI VSS TSMC_223 
+ TSMC_224 TSMC_287 TSMC_288 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO17 TSMC_29 TSMC_30 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_93 TSMC_94 TSMC_157 TSMC_158 TSMC_373 VDDM VDDAI VDDI VSS TSMC_221 
+ TSMC_222 TSMC_285 TSMC_286 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO18 TSMC_27 TSMC_28 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_91 TSMC_92 TSMC_155 TSMC_156 TSMC_373 VDDM VDDAI VDDI VSS TSMC_219 
+ TSMC_220 TSMC_283 TSMC_284 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO19 TSMC_25 TSMC_26 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_89 TSMC_90 TSMC_153 TSMC_154 TSMC_373 VDDM VDDAI VDDI VSS TSMC_217 
+ TSMC_218 TSMC_281 TSMC_282 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO20 TSMC_23 TSMC_24 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_87 TSMC_88 TSMC_151 TSMC_152 TSMC_373 VDDM VDDAI VDDI VSS TSMC_215 
+ TSMC_216 TSMC_279 TSMC_280 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO21 TSMC_21 TSMC_22 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_85 TSMC_86 TSMC_149 TSMC_150 TSMC_373 VDDM VDDAI VDDI VSS TSMC_213 
+ TSMC_214 TSMC_277 TSMC_278 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO22 TSMC_19 TSMC_20 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_83 TSMC_84 TSMC_147 TSMC_148 TSMC_373 VDDM VDDAI VDDI VSS TSMC_211 
+ TSMC_212 TSMC_275 TSMC_276 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO23 TSMC_17 TSMC_18 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_81 TSMC_82 TSMC_145 TSMC_146 TSMC_373 VDDM VDDAI VDDI VSS TSMC_209 
+ TSMC_210 TSMC_273 TSMC_274 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO24 TSMC_15 TSMC_16 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_79 TSMC_80 TSMC_143 TSMC_144 TSMC_373 VDDM VDDAI VDDI VSS TSMC_207 
+ TSMC_208 TSMC_271 TSMC_272 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO25 TSMC_13 TSMC_14 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_77 TSMC_78 TSMC_141 TSMC_142 TSMC_373 VDDM VDDAI VDDI VSS TSMC_205 
+ TSMC_206 TSMC_269 TSMC_270 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO26 TSMC_11 TSMC_12 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_75 TSMC_76 TSMC_139 TSMC_140 TSMC_373 VDDM VDDAI VDDI VSS TSMC_203 
+ TSMC_204 TSMC_267 TSMC_268 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO27 TSMC_9 TSMC_10 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_73 TSMC_74 TSMC_137 TSMC_138 TSMC_373 VDDM VDDAI VDDI VSS TSMC_201 
+ TSMC_202 TSMC_265 TSMC_266 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO28 TSMC_7 TSMC_8 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_71 TSMC_72 TSMC_135 TSMC_136 TSMC_373 VDDM VDDAI VDDI VSS TSMC_199 
+ TSMC_200 TSMC_263 TSMC_264 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO29 TSMC_5 TSMC_6 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_69 TSMC_70 TSMC_133 TSMC_134 TSMC_373 VDDM VDDAI VDDI VSS TSMC_197 
+ TSMC_198 TSMC_261 TSMC_262 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO30 TSMC_3 TSMC_4 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_67 TSMC_68 TSMC_131 TSMC_132 TSMC_373 VDDM VDDAI VDDI VSS TSMC_195 
+ TSMC_196 TSMC_259 TSMC_260 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XLIO31 TSMC_1 TSMC_2 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_65 TSMC_66 TSMC_129 TSMC_130 TSMC_373 VDDM VDDAI VDDI VSS TSMC_193 
+ TSMC_194 TSMC_257 TSMC_258 S6ALLSVTFW10V20_RF_LIOX2_72_V1 
XTROLIOL TSMC_399 TSMC_321 TSMC_397 TSMC_322 TSMC_323 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_407 TSMC_408 TSMC_409 TSMC_405 TSMC_406 TSMC_324 
+ TSMC_325 TSMC_401 TSMC_327 TSMC_373 VDDM VDDAI VDDI VSS TSMC_410 
+ TSMC_329 TSMC_411 TSMC_331 TSMC_332 TSMC_333 
+ S6ALLSVTFW10V20_RF_TRKLIOX2_72_V1 
XTROLIOR TSMC_399 TSMC_334 TSMC_412 TSMC_335 TSMC_336 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_407 TSMC_408 TSMC_409 TSMC_405 TSMC_406 TSMC_324 
+ TSMC_325 TSMC_401 TSMC_337 TSMC_373 VDDM VDDAI VDDI VSS TSMC_338 
+ TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 
+ S6ALLSVTFW10V20_RF_TRKLIOX2_72_V1 
XLCTRL TSMC_398 TSMC_344 TSMC_345 TSMC_399 TSMC_400 TSMC_413 TSMC_414 TSMC_402 
+ TSMC_403 TSMC_404 TSMC_407 TSMC_408 TSMC_409 TSMC_346 TSMC_347 
+ TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_405 TSMC_406 TSMC_324 
+ TSMC_415 TSMC_352 TSMC_326 TSMC_353 TSMC_354 TSMC_355 TSMC_356 
+ TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 TSMC_362 TSMC_363 TSMC_364 
+ TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 TSMC_370 TSMC_371 
+ TSMC_372 TSMC_373 TSMC_325 TSMC_374 TSMC_375 VDDM VDDI VSS TSMC_376 
+ TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 
+ TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 
+ TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ S6ALLSVTFW10V20_RF_LCTRL 
.ENDS

.SUBCKT S6ALLSVTFW10V20_WRITE_TRAKING TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 VDDM VDDI VDDAI VSS TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 
XRWLLD0 TSMC_63 TSMC_64 TSMC_127 TSMC_128 VSS VDDM VDDAI VSS TSMC_255 TSMC_256 
+ TSMC_191 TSMC_192 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD1 TSMC_61 TSMC_62 TSMC_125 TSMC_126 VSS VDDM VDDAI VSS TSMC_253 TSMC_254 
+ TSMC_189 TSMC_190 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD2 TSMC_59 TSMC_60 TSMC_123 TSMC_124 VSS VDDM VDDAI VSS TSMC_251 TSMC_252 
+ TSMC_187 TSMC_188 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD3 TSMC_57 TSMC_58 TSMC_121 TSMC_122 VSS VDDM VDDAI VSS TSMC_249 TSMC_250 
+ TSMC_185 TSMC_186 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD4 TSMC_55 TSMC_56 TSMC_119 TSMC_120 VSS VDDM VDDAI VSS TSMC_247 TSMC_248 
+ TSMC_183 TSMC_184 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD5 TSMC_53 TSMC_54 TSMC_117 TSMC_118 VSS VDDM VDDAI VSS TSMC_245 
+ TSMC_246 TSMC_181 TSMC_182 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD6 TSMC_51 TSMC_52 TSMC_115 TSMC_116 VSS VDDM VDDAI VSS TSMC_243 
+ TSMC_244 TSMC_179 TSMC_180 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD7 TSMC_49 TSMC_50 TSMC_113 TSMC_114 VSS VDDM VDDAI VSS TSMC_241 
+ TSMC_242 TSMC_177 TSMC_178 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD8 TSMC_47 TSMC_48 TSMC_111 TSMC_112 VSS VDDM VDDAI VSS TSMC_239 
+ TSMC_240 TSMC_175 TSMC_176 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD9 TSMC_45 TSMC_46 TSMC_109 TSMC_110 VSS VDDM VDDAI VSS TSMC_237 
+ TSMC_238 TSMC_173 TSMC_174 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD10 TSMC_43 TSMC_44 TSMC_107 TSMC_108 VSS VDDM VDDAI VSS TSMC_235 
+ TSMC_236 TSMC_171 TSMC_172 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD11 TSMC_41 TSMC_42 TSMC_105 TSMC_106 VSS VDDM VDDAI VSS TSMC_233 
+ TSMC_234 TSMC_169 TSMC_170 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD12 TSMC_39 TSMC_40 TSMC_103 TSMC_104 VSS VDDM VDDAI VSS TSMC_231 
+ TSMC_232 TSMC_167 TSMC_168 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD13 TSMC_37 TSMC_38 TSMC_101 TSMC_102 VSS VDDM VDDAI VSS TSMC_229 
+ TSMC_230 TSMC_165 TSMC_166 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD14 TSMC_35 TSMC_36 TSMC_99 TSMC_100 VSS VDDM VDDAI VSS TSMC_227 
+ TSMC_228 TSMC_163 TSMC_164 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD15 TSMC_33 TSMC_34 TSMC_97 TSMC_98 VSS VDDM VDDAI VSS TSMC_225 
+ TSMC_226 TSMC_161 TSMC_162 TSMC_273 TSMC_274 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD16 TSMC_31 TSMC_32 TSMC_95 TSMC_96 VSS VDDM VDDAI VSS TSMC_223 
+ TSMC_224 TSMC_159 TSMC_160 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD17 TSMC_29 TSMC_30 TSMC_93 TSMC_94 VSS VDDM VDDAI VSS TSMC_221 
+ TSMC_222 TSMC_157 TSMC_158 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD18 TSMC_27 TSMC_28 TSMC_91 TSMC_92 VSS VDDM VDDAI VSS TSMC_219 
+ TSMC_220 TSMC_155 TSMC_156 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD19 TSMC_25 TSMC_26 TSMC_89 TSMC_90 VSS VDDM VDDAI VSS TSMC_217 
+ TSMC_218 TSMC_153 TSMC_154 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD20 TSMC_23 TSMC_24 TSMC_87 TSMC_88 VSS VDDM VDDAI VSS TSMC_215 
+ TSMC_216 TSMC_151 TSMC_152 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD21 TSMC_21 TSMC_22 TSMC_85 TSMC_86 VSS VDDM VDDAI VSS TSMC_213 
+ TSMC_214 TSMC_149 TSMC_150 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD22 TSMC_19 TSMC_20 TSMC_83 TSMC_84 VSS VDDM VDDAI VSS TSMC_211 
+ TSMC_212 TSMC_147 TSMC_148 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD23 TSMC_17 TSMC_18 TSMC_81 TSMC_82 VSS VDDM VDDAI VSS TSMC_209 
+ TSMC_210 TSMC_145 TSMC_146 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD24 TSMC_15 TSMC_16 TSMC_79 TSMC_80 VSS VDDM VDDAI VSS TSMC_207 
+ TSMC_208 TSMC_143 TSMC_144 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD25 TSMC_13 TSMC_14 TSMC_77 TSMC_78 VSS VDDM VDDAI VSS TSMC_205 
+ TSMC_206 TSMC_141 TSMC_142 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD26 TSMC_11 TSMC_12 TSMC_75 TSMC_76 VSS VDDM VDDAI VSS TSMC_203 
+ TSMC_204 TSMC_139 TSMC_140 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD27 TSMC_9 TSMC_10 TSMC_73 TSMC_74 VSS VDDM VDDAI VSS TSMC_201 
+ TSMC_202 TSMC_137 TSMC_138 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD28 TSMC_7 TSMC_8 TSMC_71 TSMC_72 VSS VDDM VDDAI VSS TSMC_199 
+ TSMC_200 TSMC_135 TSMC_136 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD29 TSMC_5 TSMC_6 TSMC_69 TSMC_70 VSS VDDM VDDAI VSS TSMC_197 
+ TSMC_198 TSMC_133 TSMC_134 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD30 TSMC_3 TSMC_4 TSMC_67 TSMC_68 VSS VDDM VDDAI VSS TSMC_195 
+ TSMC_196 TSMC_131 TSMC_132 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLD31 TSMC_1 TSMC_2 TSMC_65 TSMC_66 VSS VDDM VDDAI VSS TSMC_193 
+ TSMC_194 TSMC_129 TSMC_130 TSMC_276 TSMC_277 TSMC_275 
+ S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X2 
XRWLLDL TSMC_257 TSMC_258 VSS VDDM VDDAI VSS TSMC_278 TSMC_259 TSMC_279 
+ TSMC_275 S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X1 
XRWLLDR TSMC_261 TSMC_258 VSS VDDM VDDAI VSS TSMC_280 TSMC_262 TSMC_279 
+ TSMC_275 S6ALLSVTFW10V20_D130_ARRAY_RWL_TRK_X1 
XDECCAP TSMC_281 TSMC_267 TSMC_264 TSMC_265 TSMC_266 VDDM VDDI VSS TSMC_259 
+ TSMC_263 TSMC_260 TSMC_268 TSMC_275 TSMC_275 
+ S6ALLSVTFW10V20_RF_XDECCAP 
.ENDS

.SUBCKT TS6N16FFCLLSVTA16X32M2FW D[31] D[30] D[29] D[28] D[27] D[26] D[25] 
+ D[24] D[23] D[22] D[21] D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] 
+ D[11] D[10] D[9] D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] Q[31] Q[30] 
+ Q[29] Q[28] Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] 
+ Q[16] Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] 
+ Q[2] Q[1] Q[0] BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] BWEB[25] 
+ BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] BWEB[18] BWEB[17] 
+ BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] BWEB[11] BWEB[10] BWEB[9] 
+ BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] BWEB[3] BWEB[2] BWEB[1] BWEB[0] AB[3] 
+ AB[2] AB[1] AB[0] CLKR REB AA[3] AA[2] AA[1] AA[0] CLKW WEB KP[2] KP[1] KP[0] 
+ WCT[1] WCT[0] RCT[1] RCT[0] VDD VSS 
XPIN_ROW D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] D[22] D[21] 
+ D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] D[10] D[9] 
+ D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] Q[31] Q[30] Q[29] Q[28] 
+ Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] Q[16] 
+ Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] 
+ Q[2] Q[1] Q[0] BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] 
+ BWEB[25] BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] 
+ BWEB[18] BWEB[17] BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] 
+ BWEB[11] BWEB[10] BWEB[9] BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] 
+ BWEB[3] BWEB[2] BWEB[1] BWEB[0] TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 AB[3] AB[2] AB[1] AB[0] CLKR REB TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 AA[3] AA[2] AA[1] AA[0] CLKW WEB KP[2] KP[1] KP[0] 
+ TSMC_1 TSMC_2 TSMC_1 RCT[1] RCT[0] WCT[1] WCT[0] TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 VSS TSMC_3 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_2 TSMC_2 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_4 
+ TSMC_5 TSMC_6 S6ALLSVTFW10V20_PIN_ROW 
XGCTRL_GIO CLKR CLKW D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] 
+ D[22] D[21] D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] 
+ D[10] D[9] D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 
+ TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 
+ TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 KP[2] KP[1] KP[0] 
+ TSMC_104 TSMC_105 TSMC_106 TSMC_1 TSMC_2 TSMC_1 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_1 Q[31] Q[30] Q[29] Q[28] Q[27] Q[26] Q[25] 
+ Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] Q[16] Q[15] Q[14] Q[13] 
+ Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] 
+ RCT[1] RCT[0] REB TSMC_112 TSMC_1 TSMC_113 TSMC_114 TSMC_115 
+ TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 AB[3] AB[2] 
+ AB[1] TSMC_1 TSMC_1 AB[0] TSMC_1 TSMC_2 TSMC_1 TSMC_132 VDD VDD VSS 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 
+ TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 
+ TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 
+ TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 
+ TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 
+ TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 WCT[1] WCT[0] 
+ WEB BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] BWEB[25] 
+ BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] BWEB[18] 
+ BWEB[17] BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] BWEB[11] 
+ BWEB[10] BWEB[9] BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] BWEB[3] BWEB[2] 
+ BWEB[1] BWEB[0] TSMC_261 TSMC_1 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 
+ TSMC_280 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 AA[3] AA[2] AA[1] TSMC_1 
+ TSMC_1 AA[0] TSMC_281 TSMC_1 TSMC_3 TSMC_282 TSMC_2 TSMC_283 TSMC_2 TSMC_2 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 
+ TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 
+ TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 
+ TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 
+ TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 TSMC_347 TSMC_1 
+ S6ALLSVTFW10V20_GCTRL_GIO 
XROW_TRACKING TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 
+ TSMC_232 TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 
+ TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 
+ TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 
+ TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 
+ TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 
+ TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 
+ TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 
+ TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 
+ TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 
+ TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 
+ TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 VDD VDD 
+ VDD VSS TSMC_112 TSMC_112 TSMC_1 TSMC_132 TSMC_348 TSMC_349 
+ S6ALLSVTFW10V20_ROW_TRACKING 
XARY4ROW_SEG0_ARY0 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
+ TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 TSMC_355 
+ TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 
+ TSMC_375 TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 
+ TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 
+ TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 
+ TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 
+ TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_133 
+ TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 
+ TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 
+ TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_414 
+ TSMC_415 TSMC_110 TSMC_103 TSMC_416 TSMC_417 TSMC_116 TSMC_117 
+ TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_1 TSMC_1 
+ VDD VDD VDD VSS TSMC_261 TSMC_262 TSMC_418 TSMC_265 TSMC_266 
+ TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 
+ TSMC_123 TSMC_127 TSMC_272 TSMC_276 TSMC_348 TSMC_419 TSMC_349 
+ TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 
+ S6ALLSVTFW10V20_ARY4ROW 
XARY4ROW_TK_SEG0_ARY1 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
+ TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 TSMC_355 
+ TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 
+ TSMC_375 TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 
+ TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 
+ TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 
+ TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 
+ TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_133 
+ TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 
+ TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 
+ TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_414 
+ TSMC_415 TSMC_110 TSMC_103 TSMC_416 TSMC_417 TSMC_116 TSMC_117 
+ TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_1 TSMC_1 
+ VDD VDD VDD VSS TSMC_261 TSMC_262 TSMC_418 TSMC_265 TSMC_266 
+ TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 
+ TSMC_122 TSMC_127 TSMC_271 TSMC_276 TSMC_419 TSMC_425 TSMC_420 
+ TSMC_426 TSMC_132 TSMC_132 TSMC_422 TSMC_427 TSMC_424 
+ TSMC_428 S6ALLSVTFW10V20_ARY4ROW_TK 
XLIO_LCTRL_SEG0 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 TSMC_355 TSMC_356 
+ TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 TSMC_362 
+ TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 
+ TSMC_382 TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 
+ TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 
+ TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 
+ TSMC_408 TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_429 
+ TSMC_430 TSMC_431 TSMC_432 TSMC_433 TSMC_434 TSMC_435 
+ TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_441 TSMC_442 
+ TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 
+ TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 
+ TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 
+ TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 
+ TSMC_488 TSMC_489 TSMC_490 TSMC_491 TSMC_492 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 
+ TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_133 TSMC_134 TSMC_135 
+ TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 
+ TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 
+ TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 
+ TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 
+ TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 
+ TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_493 TSMC_414 TSMC_493 
+ TSMC_1 TSMC_415 TSMC_112 TSMC_132 TSMC_1 TSMC_1 TSMC_1 TSMC_110 
+ TSMC_111 TSMC_132 TSMC_494 TSMC_103 TSMC_494 TSMC_132 TSMC_1 TSMC_1 
+ TSMC_1 VDD TSMC_281 TSMC_132 TSMC_127 TSMC_127 TSMC_104 TSMC_105 TSMC_106 
+ TSMC_107 TSMC_108 TSMC_109 TSMC_1 TSMC_495 TSMC_113 TSMC_417 
+ TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_1 TSMC_1 TSMC_126 TSMC_126 VDD VDD VDD VSS 
+ TSMC_261 TSMC_262 TSMC_418 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 
+ TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 
+ TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_112 TSMC_261 TSMC_496 
+ TSMC_283 TSMC_1 TSMC_497 TSMC_112 S6ALLSVTFW10V20_LIO_LCTRL 
XWRITE_TRAKING TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 TSMC_355 TSMC_356 
+ TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 TSMC_362 
+ TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 
+ TSMC_382 TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 
+ TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 
+ TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 
+ TSMC_408 TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_133 
+ TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 
+ TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 
+ TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 
+ TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 
+ TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_414 TSMC_415 
+ TSMC_110 TSMC_111 TSMC_103 TSMC_416 TSMC_281 TSMC_112 TSMC_495 
+ TSMC_1 TSMC_1 VDD VDD VDD VSS TSMC_261 TSMC_425 TSMC_426 TSMC_427 
+ TSMC_428 S6ALLSVTFW10V20_WRITE_TRAKING 
.ENDS


