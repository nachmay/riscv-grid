**** Created by MC2: Version 2013.12.00.f on 2025/06/18, 12:00:46 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  TS16FF2PRF
* Top Cell Name: all_leafcells
* View Name:     schematic
* Netlisted on:  Sep 30 16:22:09 2015
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM


*.PIN vss

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_svt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nand2_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_svt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_inv_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_svt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nor2_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WCTD VDD VDDI VSS TSMC_1 TSMC_2 TSMC_3 TSMC_4 
XI76 TSMC_5 TSMC_6 VSS VSS VDDI VDD TSMC_3 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI79 TSMC_7 TSMC_8 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI66 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_2 TSMC_11 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_7 TSMC_12 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_14 TSMC_7 VSS VSS VDDI VDD TSMC_6 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_1 TSMC_15 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_9 TSMC_16 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_17 TSMC_11 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_16 TSMC_15 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI145 VSS VSS TSMC_4 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_18 TSMC_5 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_5 TSMC_19 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_5 TSMC_20 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI143 VSS VSS TSMC_21 TSMC_22 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI159 VSS VSS TSMC_13 TSMC_23 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_22 TSMC_17 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_24 TSMC_25 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI89 VSS VSS TSMC_10 TSMC_12 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI160 VSS VSS TSMC_13 TSMC_24 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI144 VSS VSS TSMC_25 TSMC_21 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW40W20_nor2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WRTRKEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WRTRKEN TSMC_1 VDD VDDI VSS TSMC_2 TSMC_3 TSMC_4 
XI19<0> TSMC_2 TSMC_5 VSS VSS VDDI VDD TSMC_1 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI19<1> TSMC_2 TSMC_5 VSS VSS VDDI VDD TSMC_1 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI14 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_5 
+ S6ALLSVTFW40W20_nor2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_W1TRKWR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_W1TRKWR TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS TSMC_4 
+ TSMC_5 
XXwctd VDD VDDI VSS TSMC_1 TSMC_2 TSMC_6 TSMC_4 S6ALLSVTFW40W20_RF_WCTD 
XXrdtrken TSMC_3 VDD VDDI VSS TSMC_6 TSMC_4 TSMC_5 
+ S6ALLSVTFW40W20_RF_WRTRKEN 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WREFMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WREFMUX TSMC_1 VDD VDDI VSS TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
MM10 TSMC_7 TSMC_1 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_4 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_4 TSMC_6 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM13 TSMC_8 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_3 TSMC_6 TSMC_9 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM12 TSMC_9 TSMC_1 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_3 TSMC_5 TSMC_4 VDD pch_svt_mac l=0.020u nfin=3 m=2 
MM9 TSMC_3 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM8 TSMC_4 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM0 TSMC_3 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_1 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_3 TSMC_10 TSMC_2 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM5 TSMC_4 TSMC_11 TSMC_2 VSS nch_svt_mac l=0.020u nfin=6 m=2 
XI21 TSMC_6 TSMC_7 TSMC_2 VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI19 TSMC_6 TSMC_1 TSMC_2 VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKGIOWR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TRKGIOWR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 
XXwrst TSMC_15 TSMC_16 TSMC_20 VDD VDDI VSS TSMC_17 TSMC_29 
+ S6ALLSVTFW40W20_RF_W1TRKWR 
XXwrefmux TSMC_11 VDD VDDI VSS VSS TSMC_12 TSMC_14 TSMC_30 TSMC_29 
+ S6ALLSVTFW40W20_RF_WREFMUX 
XI21 VSS VSS TSMC_19 TSMC_29 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_29 TSMC_30 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 p_nfin=7 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WMUX TSMC_1 TSMC_2 VDD VDDI VSS TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM0 TSMC_4 TSMC_8 TSMC_3 VSS nch_lvt_mac l=0.020u nfin=6 m=2 
MM2 TSMC_5 TSMC_9 TSMC_3 VSS nch_lvt_mac l=0.020u nfin=6 m=2 
MM13 TSMC_10 TSMC_1 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_4 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_4 TSMC_11 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_5 TSMC_11 TSMC_10 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM9 TSMC_4 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM4 TSMC_5 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM10 TSMC_4 TSMC_6 TSMC_5 VDD pch_svt_mac l=0.020u nfin=3 m=2 
MM6 TSMC_5 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM12 TSMC_12 TSMC_2 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI23 VSS VSS TSMC_7 TSMC_11 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI14 TSMC_11 TSMC_2 TSMC_3 VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI15 TSMC_11 TSMC_1 TSMC_3 VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRI_W3L2M1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TRI_W3L2M1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM4 TSMC_9 TSMC_7 TSMC_4 TSMC_5 pch_svt_mac l=0.020u nfin=3 m=1 
MM5 TSMC_8 TSMC_1 TSMC_9 TSMC_5 pch_svt_mac l=0.020u nfin=3 m=1 
MM6 TSMC_10 TSMC_6 TSMC_2 TSMC_3 nch_svt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_8 TSMC_1 TSMC_10 TSMC_3 nch_svt_mac l=0.020u nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRI_W2L2M1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TRI_W2L2M1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM4 TSMC_9 TSMC_7 TSMC_4 TSMC_5 pch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_8 TSMC_1 TSMC_9 TSMC_5 pch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_10 TSMC_6 TSMC_2 TSMC_3 nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_8 TSMC_1 TSMC_10 TSMC_3 nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DIN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_DIN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD 
+ VDDI VSS TSMC_7 
XI16 TSMC_8 VSS VSS VDDI VDD TSMC_4 TSMC_5 TSMC_9 
+ S6ALLSVTFW40W20_RF_TRI_W3L2M1 
XI90 TSMC_10 VSS VSS VDDI VDD TSMC_4 TSMC_5 TSMC_11 
+ S6ALLSVTFW40W20_RF_TRI_W3L2M1 
XI15 TSMC_12 TSMC_13 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_12 TSMC_14 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI63 VSS VSS TSMC_15 TSMC_12 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI59 VSS VSS TSMC_16 TSMC_14 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI61 VSS VSS TSMC_7 TSMC_17 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI83 VSS VSS TSMC_9 TSMC_3 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI92 VSS VSS TSMC_11 TSMC_2 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI99 VSS VSS TSMC_1 TSMC_16 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI62 VSS VSS TSMC_17 TSMC_15 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI60 VSS VSS TSMC_14 TSMC_13 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI94 TSMC_2 VSS VSS VDDI VDD TSMC_5 TSMC_4 TSMC_11 
+ S6ALLSVTFW40W20_RF_TRI_W2L2M1 
XI17 TSMC_3 VSS VSS VDDI VDD TSMC_5 TSMC_4 TSMC_9 
+ S6ALLSVTFW40W20_RF_TRI_W2L2M1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DOLATCHM48
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_DOLATCHM48 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 
MM0 TSMC_3 TSMC_4 VDD VDD pch_svt_mac l=0.020u nfin=3 m=1 
XI3 VSS VSS TSMC_3 TSMC_1 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI7 TSMC_2 VSS VSS VDDI VDD TSMC_5 TSMC_6 TSMC_3 
+ S6ALLSVTFW40W20_RF_TRI_W3L2M1 
XI5 TSMC_3 VSS VSS VDDI VDD TSMC_7 TSMC_8 TSMC_2 
+ S6ALLSVTFW40W20_RF_TRI_W3L2M1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DINM4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_DINM4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
XI19 VSS VSS TSMC_18 TSMC_24 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI20 VSS VSS TSMC_24 TSMC_25 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI18<1> VSS VSS TSMC_19 TSMC_26 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI18<0> VSS VSS TSMC_19 TSMC_27 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI15<1> VSS VSS TSMC_26 TSMC_28 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=7 p_l=0.020u 
XI15<0> VSS VSS TSMC_27 TSMC_29 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=7 p_l=0.020u 
XXdltch TSMC_1 TSMC_2 TSMC_3 TSMC_24 TSMC_25 TSMC_4 VDD VDDI VSS TSMC_17 
+ S6ALLSVTFW40W20_RF_DIN 
XXwmux<2> TSMC_2 TSMC_3 VDD VDDI VSS TSMC_6 TSMC_10 TSMC_14 TSMC_28 
+ TSMC_21 S6ALLSVTFW40W20_RF_WMUX 
XXwmux<1> TSMC_2 TSMC_3 VDD VDDI VSS TSMC_7 TSMC_11 TSMC_15 TSMC_29 
+ TSMC_22 S6ALLSVTFW40W20_RF_WMUX 
XXwmux<0> TSMC_2 TSMC_3 VDD VDDI VSS TSMC_8 TSMC_12 TSMC_16 TSMC_29 
+ TSMC_23 S6ALLSVTFW40W20_RF_WMUX 
XXwmux_f TSMC_2 TSMC_3 VDD VDDI VSS TSMC_5 TSMC_9 TSMC_13 TSMC_28 
+ TSMC_20 S6ALLSVTFW40W20_RF_WMUX 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    TRI_M4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_TRI_M4 TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS TSMC_4 
MM3 TSMC_4 TSMC_3 TSMC_5 VDD pch_lvt_mac l=0.020u nfin=4 m=3 
MM0 TSMC_5 TSMC_1 VDDI VDD pch_lvt_mac l=0.020u nfin=4 m=3 
MM1 TSMC_4 TSMC_2 TSMC_6 VSS nch_svt_mac l=0.020u nfin=4 m=2 
MM2 TSMC_6 TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=4 m=2 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RMUX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RMUX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
XI9 TSMC_1 TSMC_5 TSMC_4 VDD VDDI VSS TSMC_2 S6ALLSVTFW40W20_TRI_M4 
MM1 TSMC_1 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=4 m=3 
MM5 TSMC_6 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_1 TSMC_7 TSMC_6 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI1 VSS VSS TSMC_1 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
MM2 TSMC_1 TSMC_7 TSMC_8 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_8 TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DOUTM4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_DOUTM4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDI VSS TSMC_13 TSMC_14 
MM4 TSMC_15 TSMC_16 VDD VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_15 TSMC_6 VDD VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_16 TSMC_12 VDD VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_16 TSMC_13 VDD VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_15 TSMC_6 TSMC_17 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_16 TSMC_13 TSMC_18 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_18 TSMC_12 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_17 TSMC_16 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
XXrmux<2> TSMC_3 TSMC_19 TSMC_20 TSMC_21 TSMC_22 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_RMUX4 
XXrmux<1> TSMC_4 TSMC_19 TSMC_20 TSMC_23 TSMC_24 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_RMUX4 
XXrmux<0> TSMC_5 TSMC_19 TSMC_20 TSMC_25 TSMC_26 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_RMUX4 
XXrmux_f TSMC_2 TSMC_19 TSMC_20 TSMC_27 TSMC_28 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_RMUX4 
XXqltch TSMC_7 TSMC_1 TSMC_19 TSMC_6 TSMC_29 TSMC_15 VDD VDDI VSS TSMC_13 
+ TSMC_14 S6ALLSVTFW40W20_RF_DOLATCHM48 
XI27<3> VSS VSS TSMC_28 TSMC_27 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI27<2> VSS VSS TSMC_22 TSMC_21 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI27<1> VSS VSS TSMC_24 TSMC_23 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI27<0> VSS VSS TSMC_26 TSMC_25 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI10 VSS VSS TSMC_15 TSMC_30 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI13 VSS VSS TSMC_15 TSMC_29 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI29 VSS VSS TSMC_30 TSMC_20 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=5 p_l=0.020u 
XI28<3> TSMC_8 TSMC_16 VSS VSS VDD VDD TSMC_28 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI28<2> TSMC_9 TSMC_16 VSS VSS VDD VDD TSMC_22 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI28<1> TSMC_10 TSMC_16 VSS VSS VDD VDD TSMC_24 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI28<0> TSMC_11 TSMC_16 VSS VSS VDD VDD TSMC_26 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_GIOM4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_GIOM4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ VDD VDDI VSS TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 
XXdin TSMC_1 TSMC_7 TSMC_8 TSMC_16 VDD VDDI VSS TSMC_17 TSMC_17 TSMC_17 TSMC_17 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 
+ TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ S6ALLSVTFW40W20_RF_DINM4 
XXdout TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_35 TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 TSMC_14 TSMC_15 VDD VDDI VSS TSMC_18 TSMC_19 
+ S6ALLSVTFW40W20_RF_DOUTM4 
XI26 VSS VSS TSMC_9 TSMC_35 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_svt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nand3_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RLCTRL_DK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RLCTRL_DK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 VDD VDDI VSS TSMC_27 
MM12 TSMC_28 TSMC_29 TSMC_30 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM11 TSMC_30 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM7 TSMC_32 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM6 TSMC_33 TSMC_34 TSMC_32 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM5 TSMC_33 TSMC_35 TSMC_32 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM1 TSMC_36 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=8 m=16 
MM0 TSMC_36 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=8 m=16 
MM8 TSMC_28 TSMC_35 TSMC_30 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM13 TSMC_28 TSMC_31 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM4 TSMC_33 TSMC_31 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM3 TSMC_33 TSMC_35 TSMC_37 VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM2 TSMC_37 TSMC_34 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM10 TSMC_38 TSMC_29 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM9 TSMC_28 TSMC_35 TSMC_38 VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
XI96 TSMC_36 VSS TSMC_39 TSMC_18 VDD VDD 
+ S6ALLSVTFW40W20_inv_ulvt_mac_pcell n_totalM=16 n_nfin=6 n_l=0.020u 
+ p_totalM=16 p_nfin=6 p_l=0.020u 
XI100 VSS VSS TSMC_1 TSMC_40 VDDI VDD 
+ S6ALLSVTFW40W20_inv_ulvt_mac_pcell n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI107 VSS VSS TSMC_41 TSMC_5 VDD VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI91 VSS VSS TSMC_33 TSMC_42 VDD VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=5 n_nfin=7 n_l=0.020u p_totalM=5 p_nfin=6 p_l=0.020u 
XI92 TSMC_36 VSS TSMC_42 TSMC_19 VDD VDD 
+ S6ALLSVTFW40W20_inv_ulvt_mac_pcell n_totalM=16 n_nfin=6 n_l=0.020u 
+ p_totalM=16 p_nfin=6 p_l=0.020u 
XI106 VSS VSS TSMC_4 TSMC_41 VDD VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI98 VSS VSS TSMC_35 TSMC_23 VDDI VDD 
+ S6ALLSVTFW40W20_inv_ulvt_mac_pcell n_totalM=14 n_nfin=5 n_l=0.020u 
+ p_totalM=14 p_nfin=5 p_l=0.020u 
XI101 VSS VSS TSMC_40 TSMC_11 VDDI VDD 
+ S6ALLSVTFW40W20_inv_ulvt_mac_pcell n_totalM=10 n_nfin=7 n_l=0.020u 
+ p_totalM=10 p_nfin=8 p_l=0.020u 
XI93_Lg16 TSMC_21 TSMC_22 TSMC_27 VSS VSS VDD VDD TSMC_35 
+ S6ALLSVTFW40W20_nand3_ulvt_mac_pcell n_totalM=4 n_nfin=7 n_l=0.020u 
+ p_totalM=4 p_nfin=2 p_l=0.020u 
XI95 TSMC_25 TSMC_26 VSS VSS VDDI VDD TSMC_34 
+ S6ALLSVTFW40W20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI103 TSMC_28 TSMC_24 VSS VSS VDD VDD TSMC_39 
+ S6ALLSVTFW40W20_nor2_ulvt_mac_pcell n_totalM=6 n_nfin=6 n_l=0.020u p_totalM=6 
+ p_nfin=7 p_l=0.020u 
XI102 TSMC_4 TSMC_4 VSS VSS VDD VDD TSMC_31 
+ S6ALLSVTFW40W20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI99 TSMC_2 TSMC_3 VSS VSS VDDI VDD TSMC_29 
+ S6ALLSVTFW40W20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WLCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WLCTRL VDD VDDI VSS TSMC_1 TSMC_2 TSMC_3 TSMC_4 
XI27 TSMC_1 TSMC_2 TSMC_4 VSS VSS VDD VDD TSMC_5 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=4 n_nfin=7 n_l=0.020u p_totalM=4 
+ p_nfin=2 p_l=0.020u 
XI28 VSS VSS TSMC_5 TSMC_3 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=14 n_nfin=5 n_l=0.020u p_totalM=14 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LCTRL_DK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_LCTRL_DK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
MM6 TSMC_71 TSMC_46 VDD VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM4 VDDI TSMC_46 VDDI VDD pch_ulvt_mac l=0.020u nfin=8 m=2 
MM5 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=12 m=16 
MM1 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=5 m=16 
MM0 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=9 m=32 
MM2 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=10 m=16 
XXrlctrl TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_17 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_25 TSMC_27 TSMC_28 TSMC_45 TSMC_48 TSMC_49 VDD 
+ VDDI VSS TSMC_69 S6ALLSVTFW40W20_RF_RLCTRL_DK 
XXwlctrl VDD VDDI VSS TSMC_50 TSMC_51 TSMC_52 TSMC_70 
+ S6ALLSVTFW40W20_RF_WLCTRL 
XI51 VSS VSS TSMC_73 TSMC_72 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI52 TSMC_24 TSMC_4 VSS VSS VDD VDD TSMC_73 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
MM3 VSS TSMC_46 VSS VSS nch_ulvt_mac l=0.020u nfin=7 m=2 
MM7 TSMC_46 TSMC_71 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_LCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
XI152 TSMC_15 TSMC_24 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=2 n_nfin=12 n_l=0.020u p_totalM=2 
+ p_nfin=12 p_l=0.020u 
XI49<1> VSS VSS TSMC_18 TSMC_12 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI49<0> VSS VSS TSMC_19 TSMC_13 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
Xlctrl TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ S6ALLSVTFW40W20_RF_LCTRL_DK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_XDECCAP
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_XDECCAP TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 
MM0_LVT TSMC_12 TSMC_6 VSS VSS nch_lvt_mac l=0.020u nfin=5 m=1 
MM196_LVT TSMC_13 TSMC_12 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM197_LVT TSMC_14 TSMC_12 TSMC_13 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM194_LVT TSMC_12 TSMC_15 VSS VSS nch_lvt_mac l=0.020u nfin=5 m=1 
MM4 TSMC_10 TSMC_16 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MMWLDRPCHWTK TSMC_10 TSMC_16 VDDI VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM195_LVT TSMC_14 TSMC_12 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=2 
MM198_LVT TSMC_17 TSMC_15 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM193_LVT TSMC_12 TSMC_6 TSMC_17 VDD pch_lvt_mac l=0.020u nfin=2 m=1 
XI78 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=6 n_l=0.020u p_totalM=2 p_nfin=6 p_l=0.020u 
XI75 VSS VSS TSMC_9 TSMC_18 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI79 VSS VSS TSMC_3 TSMC_4 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI72_LVT VSS VSS TSMC_11 TSMC_15 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI73_LVT VSS VSS TSMC_14 TSMC_19 VDDI VDD 
+ S6ALLSVTFW40W20_inv_lvt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI77 VSS VSS TSMC_2 TSMC_20 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI76 VSS VSS TSMC_18 TSMC_21 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI81_LVT TSMC_10 TSMC_19 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=8 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI82 TSMC_20 TSMC_21 VSS VSS VDD VDD TSMC_16 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=12 n_l=0.020u 
+ p_totalM=1 p_nfin=10 p_l=0.020u 
XI80_LVT TSMC_10 TSMC_19 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=6 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TRKCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 VDD VDDI VSS TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 
MM4 TSMC_37 TSMC_56 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
XI76 VSS VSS TSMC_57 TSMC_58 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI75 VSS VSS TSMC_12 TSMC_57 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI78 TSMC_13 TSMC_14 VSS VSS VDD VDD TSMC_56 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=12 n_l=0.020u 
+ p_totalM=1 p_nfin=6 p_l=0.020u 
XI79 TSMC_58 TSMC_14 VSS VSS VDDI VDD TSMC_59 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=7 p_l=0.020u 
MMWLDRPCHRTK TSMC_37 TSMC_56 VDDI VDD pch_svt_mac l=0.020u nfin=11 m=4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WXDEC TSMC_1 TSMC_2 TSMC_3 VDD VDDI TSMC_4 VSS 
+ TSMC_5 TSMC_6 
MM3 TSMC_1 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM2 TSMC_7 TSMC_8 TSMC_1 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM4 TSMC_5 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MMWLDRPCH TSMC_5 TSMC_7 TSMC_4 VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MM0 TSMC_7 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
XI58<1> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI58<0> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDECX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WXDECX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XI64<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XIXDEC<3> TSMC_16 TSMC_2 TSMC_3 VDD VDDI TSMC_7 VSS TSMC_8 TSMC_15 
+ S6ALLSVTFW40W20_RF_WXDEC 
XIXDEC<1> TSMC_16 TSMC_2 TSMC_5 VDD VDDI TSMC_7 VSS TSMC_10 TSMC_15 
+ S6ALLSVTFW40W20_RF_WXDEC 
XIXDEC<0> TSMC_17 TSMC_1 TSMC_6 VDD VDDI TSMC_7 VSS TSMC_11 TSMC_14 
+ S6ALLSVTFW40W20_RF_WXDEC 
XIXDEC<2> TSMC_17 TSMC_1 TSMC_4 VDD VDDI TSMC_7 VSS TSMC_9 TSMC_14 
+ S6ALLSVTFW40W20_RF_WXDEC 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDECX4_LR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WXDECX4_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD VDDI TSMC_7 VSS 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ S6ALLSVTFW40W20_RF_WXDECX4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RXDEC TSMC_1 TSMC_2 TSMC_3 VDD VDDI TSMC_4 VSS 
+ TSMC_5 TSMC_6 
MM1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MMWLDRPCH TSMC_5 TSMC_7 TSMC_4 VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM0 TSMC_7 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MM4 TSMC_5 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MM2 TSMC_7 TSMC_8 TSMC_1 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM3 TSMC_1 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=6 m=2 
XI58<1> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI58<0> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDECX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RXDECX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC<1> TSMC_14 TSMC_2 TSMC_5 VDD VDDI TSMC_7 VSS TSMC_10 TSMC_15 
+ S6ALLSVTFW40W20_RF_RXDEC 
XIXDEC<3> TSMC_14 TSMC_2 TSMC_3 VDD VDDI TSMC_7 VSS TSMC_8 TSMC_15 
+ S6ALLSVTFW40W20_RF_RXDEC 
XIXDEC<2> TSMC_16 TSMC_1 TSMC_4 VDD VDDI TSMC_7 VSS TSMC_9 TSMC_17 
+ S6ALLSVTFW40W20_RF_RXDEC 
XIXDEC<0> TSMC_16 TSMC_1 TSMC_6 VDD VDDI TSMC_7 VSS TSMC_11 TSMC_17 
+ S6ALLSVTFW40W20_RF_RXDEC 
XI64<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDECX4_LR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RXDECX4_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD VDDI TSMC_7 VSS 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ S6ALLSVTFW40W20_RF_RXDECX4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_XDEC4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_XDEC4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 VDD VDDI TSMC_42 VSS 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
XXwdec TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 VDD VDDI TSMC_42 VSS 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_69 TSMC_70 
+ S6ALLSVTFW40W20_RF_WXDECX4_LR 
XXrdec TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 VDD VDDI TSMC_42 VSS 
+ TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_67 TSMC_68 
+ S6ALLSVTFW40W20_RF_RXDECX4_LR 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TIELGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TIELGEN TSMC_1 TSMC_2 VDD VSS 
MM5 TSMC_1 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_3 TSMC_4 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_2 TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=3 m=2 
MM2 TSMC_3 TSMC_5 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_2 TSMC_6 VSS VSS nch_svt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_3 TSMC_5 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI0 VSS VSS TSMC_5 TSMC_4 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI1 VSS VSS TSMC_4 TSMC_6 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PUDELAY
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_PUDELAY TSMC_1 TSMC_2 TSMC_3 VDD VSS 
XI3 VSS VSS TSMC_4 TSMC_2 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI149 TSMC_1 TSMC_3 VSS VSS VDD VDD TSMC_4 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DEC2TO4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_DEC2TO4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS 
XI26 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI27 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI28 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI33 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI34 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI37 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI31 VSS VSS TSMC_10 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI35 VSS VSS TSMC_11 TSMC_6 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI39 VSS VSS TSMC_12 TSMC_5 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI29 VSS VSS TSMC_9 TSMC_8 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_YDEC3TO8L
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_YDEC3TO8L TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
XI32 TSMC_3 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI42 TSMC_6 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI38 TSMC_6 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI43 TSMC_3 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI39 TSMC_3 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_19 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI35 TSMC_6 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_3 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_6 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 VSS VSS TSMC_17 TSMC_23 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI82 VSS VSS TSMC_24 TSMC_12 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI15 VSS VSS TSMC_25 TSMC_14 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI85 VSS VSS TSMC_26 TSMC_9 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI3 VSS VSS TSMC_22 TSMC_25 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI94 VSS VSS TSMC_18 TSMC_27 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI93 VSS VSS TSMC_16 TSMC_28 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI81 VSS VSS TSMC_29 TSMC_13 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI87 VSS VSS TSMC_27 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI92 VSS VSS TSMC_19 TSMC_26 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI90 VSS VSS TSMC_21 TSMC_30 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI83 VSS VSS TSMC_30 TSMC_11 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI84 VSS VSS TSMC_23 TSMC_10 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI89 VSS VSS TSMC_20 TSMC_24 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI88 VSS VSS TSMC_15 TSMC_29 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI86 VSS VSS TSMC_28 TSMC_8 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DECPDA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_DECPDA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS 
XI58 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI60 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI59 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI61 VSS VSS TSMC_9 TSMC_13 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI64 VSS VSS TSMC_11 TSMC_14 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI66 VSS VSS TSMC_15 TSMC_5 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI62 VSS VSS TSMC_13 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI63 VSS VSS TSMC_14 TSMC_6 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI65 VSS VSS TSMC_10 TSMC_15 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI35 VSS VSS TSMC_16 TSMC_8 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI42 VSS VSS TSMC_12 TSMC_16 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RPREDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RPREDEC TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI VSS TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 
XXpb TSMC_5 TSMC_6 TSMC_13 TSMC_14 TSMC_27 TSMC_28 TSMC_29 TSMC_30 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DEC2TO4 
XXpd TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DEC2TO4 
XXpc TSMC_3 TSMC_4 TSMC_11 TSMC_12 TSMC_31 TSMC_32 TSMC_33 TSMC_34 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DEC2TO4 
XXya TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 VDD VDDI VSS TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ S6ALLSVTFW40W20_RF_YDEC3TO8L 
XXpa TSMC_7 TSMC_8 TSMC_15 TSMC_16 TSMC_23 TSMC_24 TSMC_25 TSMC_26 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DECPDA 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RPRCHBUF
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RPRCHBUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_1 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI43 VSS VSS TSMC_3 TSMC_7 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=6 n_l=0.020u p_totalM=3 p_nfin=4 p_l=0.020u 
XI42 VSS VSS TSMC_1 TSMC_2 TSMC_6 VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI2 VSS VSS TSMC_7 TSMC_4 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=13 n_nfin=5 n_l=0.020u p_totalM=13 p_nfin=9 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RCLKGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RCLKGEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS 
XI53 TSMC_11 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW40W20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=8 p_l=0.016u 
XI25 TSMC_13 TSMC_2 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
XI73 VSS VSS TSMC_9 TSMC_15 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI5 VSS VSS TSMC_13 TSMC_16 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI6 VSS VSS TSMC_13 TSMC_3 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=9 n_nfin=5 n_l=0.016u p_totalM=9 p_nfin=5 p_l=0.016u 
XI40 VSS VSS TSMC_12 TSMC_17 VDDI VDD 
+ S6ALLSVTFW40W20_inv_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI2 VSS VSS TSMC_18 TSMC_19 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI29 VSS VSS TSMC_2 TSMC_20 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI19 VSS VSS TSMC_1 TSMC_2 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI79 VSS VSS TSMC_7 TSMC_6 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=2 n_nfin=5 n_l=0.016u p_totalM=2 p_nfin=5 p_l=0.016u 
XI17 VSS VSS TSMC_15 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=2 n_nfin=8 n_l=0.016u p_totalM=2 p_nfin=8 p_l=0.016u 
MM1 TSMC_21 TSMC_22 VDD VDD pch_ulvt_mac l=0.016u nfin=8 m=3 
MM3 TSMC_13 TSMC_4 TSMC_21 VDD pch_ulvt_mac l=0.016u nfin=8 m=3 
MM9 TSMC_18 TSMC_8 TSMC_23 VDD pch_ulvt_mac l=0.016u nfin=6 m=1 
MM5 TSMC_23 TSMC_20 VDDI VDD pch_ulvt_mac l=0.016u nfin=6 m=1 
MM13 TSMC_24 TSMC_12 VDD VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM6 TSMC_18 TSMC_19 TSMC_25 VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM12 TSMC_13 TSMC_16 TSMC_24 VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM10 TSMC_25 TSMC_14 VDDI VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM0 TSMC_16 TSMC_8 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=2 
MM8 TSMC_13 TSMC_12 VSS VSS nch_ulvt_mac l=0.016u nfin=5 m=6 
MM4 TSMC_26 TSMC_20 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM11 TSMC_18 TSMC_8 VSS VSS nch_ulvt_mac l=0.016u nfin=4 m=1 
MM2 TSMC_18 TSMC_14 VSS VSS nch_ulvt_mac l=0.016u nfin=4 m=1 
MM15 TSMC_27 TSMC_16 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM7 TSMC_18 TSMC_19 TSMC_26 VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM14 TSMC_13 TSMC_16 TSMC_27 VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
XI71 TSMC_13 TSMC_28 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nand2_ulvt_mac_pcell n_totalM=2 n_nfin=3 n_l=0.016u 
+ p_totalM=2 p_nfin=3 p_l=0.016u 
XI75 TSMC_5 TSMC_20 VSS VSS VDD VDD TSMC_28 
+ S6ALLSVTFW40W20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u 
+ p_totalM=1 p_nfin=2 p_l=0.016u 
XI56 TSMC_18 TSMC_5 VSS VSS VDD VDD TSMC_11 
+ S6ALLSVTFW40W20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u 
+ p_totalM=1 p_nfin=2 p_l=0.016u 
XI82 TSMC_29 TSMC_17 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW40W20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u 
+ p_totalM=1 p_nfin=3 p_l=0.016u 
XI8 TSMC_20 TSMC_10 VSS VSS VDDI VDD TSMC_29 
+ S6ALLSVTFW40W20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u 
+ p_totalM=1 p_nfin=2 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH_RA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_ILATCH_RA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_ulvt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_ulvt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW40W20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_ulvt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_ulvt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH_RA_Y
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_ILATCH_RA_Y TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_lvt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_lvt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW40W20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_lvt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_lvt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ADRLAT_RA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_ADRLAT_RA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 VDD VDDI VSS 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 
XXxlat<7> TSMC_25 TSMC_1 TSMC_2 TSMC_3 TSMC_11 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXxlat<6> TSMC_26 TSMC_1 TSMC_2 TSMC_4 TSMC_12 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXxlat<5> TSMC_27 TSMC_1 TSMC_2 TSMC_5 TSMC_13 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXxlat<4> TSMC_28 TSMC_1 TSMC_2 TSMC_6 TSMC_14 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXxlat<3> TSMC_29 TSMC_1 TSMC_2 TSMC_7 TSMC_15 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXxlat<2> TSMC_30 TSMC_1 TSMC_2 TSMC_8 TSMC_16 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXxlat<1> TSMC_31 TSMC_1 TSMC_2 TSMC_9 TSMC_17 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXxlat<0> TSMC_32 TSMC_1 TSMC_2 TSMC_10 TSMC_18 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA 
XXylat<2> TSMC_33 TSMC_1 TSMC_2 TSMC_19 TSMC_22 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA_Y 
XXylat<1> TSMC_34 TSMC_1 TSMC_2 TSMC_20 TSMC_23 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA_Y 
XXylat<0> TSMC_35 TSMC_1 TSMC_2 TSMC_21 TSMC_24 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH_RA_Y 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RENLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RENLAT TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
XI15 VSS VSS TSMC_5 TSMC_3 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI0 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI5 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
MM4 TSMC_8 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_9 TSMC_5 TSMC_8 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_10 TSMC_6 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_9 TSMC_2 TSMC_10 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_9 TSMC_5 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_11 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_9 TSMC_2 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_12 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI6 TSMC_4 TSMC_9 VSS VSS VDD VDD TSMC_5 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RTUNE
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RTUNE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDI VSS 
XXenlat TSMC_1 TSMC_10 TSMC_8 TSMC_9 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_RENLAT 
XI12<2> VSS VSS TSMC_13 TSMC_5 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI12<1> VSS VSS TSMC_14 TSMC_6 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI12<0> VSS VSS TSMC_15 TSMC_7 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI13<2> VSS VSS TSMC_2 TSMC_13 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI13<1> VSS VSS TSMC_3 TSMC_14 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI13<0> VSS VSS TSMC_4 TSMC_15 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI7 VSS VSS TSMC_11 TSMC_12 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=5 n_l=0.020u p_totalM=4 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RGCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RGCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 VDD VDDI VSS TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
XXpredecs TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
+ TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 VDD VDDI VSS TSMC_58 
+ TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ S6ALLSVTFW40W20_RF_RPREDEC 
XXrprchb TSMC_38 TSMC_82 TSMC_83 TSMC_43 TSMC_46 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_RPRCHBUF 
XXclkgen TSMC_1 TSMC_84 TSMC_40 TSMC_44 TSMC_85 TSMC_8 TSMC_9 TSMC_38 TSMC_83 
+ TSMC_45 VDD VDDI VSS S6ALLSVTFW40W20_RF_RCLKGEN 
XXadrlat TSMC_8 TSMC_9 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 VDD VDDI VSS 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 S6ALLSVTFW40W20_RF_ADRLAT_RA 
XXrtune TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_85 
+ TSMC_82 TSMC_39 TSMC_41 TSMC_42 VDD VDDI VSS S6ALLSVTFW40W20_RF_RTUNE 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DKCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_DKCTD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM2 VDDI TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=4 m=1 
MM1 VSS TSMC_5 VSS VSS nch_svt_mac l=0.020u nfin=4 m=1 
XI126 TSMC_4 TSMC_5 VSS VSS VDDI VDD TSMC_6 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI64 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_7 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI76 TSMC_8 TSMC_9 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI66 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_12 TSMC_6 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI179 TSMC_14 TSMC_6 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI178 TSMC_16 TSMC_6 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_1 TSMC_18 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_2 TSMC_19 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI156 TSMC_6 TSMC_10 VSS VSS VDDI VDD TSMC_3 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=6 n_nfin=10 n_l=0.020u 
+ p_totalM=6 p_nfin=5 p_l=0.020u 
XI89 VSS VSS TSMC_11 TSMC_12 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_7 TSMC_8 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_15 TSMC_20 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_21 TSMC_19 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_17 TSMC_22 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_20 TSMC_18 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_22 TSMC_9 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_13 TSMC_21 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WCLKGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WCLKGEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS TSMC_9 
MM11 TSMC_10 TSMC_11 TSMC_12 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM10 TSMC_12 TSMC_13 VDDI VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM13 TSMC_14 TSMC_15 VDD VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM2 TSMC_16 TSMC_17 VDDI VDD pch_svt_mac l=0.016u nfin=6 m=1 
MM3 TSMC_18 TSMC_3 TSMC_19 VDD pch_svt_mac l=0.016u nfin=8 m=3 
MM1 TSMC_19 TSMC_20 VDD VDD pch_svt_mac l=0.016u nfin=8 m=3 
MM0 TSMC_10 TSMC_7 TSMC_16 VDD pch_svt_mac l=0.016u nfin=6 m=1 
MM12 TSMC_18 TSMC_21 TSMC_14 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM15 TSMC_22 TSMC_21 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM7 TSMC_10 TSMC_11 TSMC_23 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM14 TSMC_18 TSMC_21 TSMC_22 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM4 TSMC_23 TSMC_17 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM9 TSMC_21 TSMC_7 VSS VSS nch_svt_mac l=0.016u nfin=2 m=2 
MM8 TSMC_18 TSMC_15 VSS VSS nch_svt_mac l=0.016u nfin=5 m=6 
MM5 TSMC_10 TSMC_7 VSS VSS nch_svt_mac l=0.016u nfin=4 m=1 
MM6 TSMC_10 TSMC_13 VSS VSS nch_svt_mac l=0.016u nfin=4 m=1 
XI61 VSS VSS TSMC_24 TSMC_9 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=5 n_l=0.016u p_totalM=6 p_nfin=5 p_l=0.016u 
XI48 VSS VSS TSMC_18 TSMC_6 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=8 n_l=0.016u p_totalM=3 p_nfin=9 p_l=0.016u 
XI45 VSS VSS TSMC_18 TSMC_25 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI28 VSS VSS TSMC_26 TSMC_24 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=8 n_l=0.016u p_totalM=1 p_nfin=8 p_l=0.016u 
XI17 VSS VSS TSMC_6 TSMC_5 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=8 n_l=0.016u p_totalM=1 p_nfin=8 p_l=0.016u 
XI44 VSS VSS TSMC_25 TSMC_27 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.016u p_totalM=2 p_nfin=4 p_l=0.016u 
XI5 VSS VSS TSMC_18 TSMC_21 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI29 VSS VSS TSMC_18 TSMC_26 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI6 VSS VSS TSMC_27 TSMC_2 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=5 n_l=0.016u p_totalM=6 p_nfin=5 p_l=0.016u 
XI26 VSS VSS TSMC_24 TSMC_9 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.016u p_totalM=4 p_nfin=8 p_l=0.016u 
XI2 VSS VSS TSMC_10 TSMC_11 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI1 VSS VSS TSMC_28 TSMC_17 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI0 VSS VSS TSMC_1 TSMC_28 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI40 VSS VSS TSMC_15 TSMC_29 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI8 TSMC_17 TSMC_8 VSS VSS VDDI VDD TSMC_30 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI37 TSMC_30 TSMC_29 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
XI52 TSMC_10 TSMC_4 VSS VSS VDD VDD TSMC_31 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI53 TSMC_31 TSMC_28 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=8 p_l=0.016u 
XI50 TSMC_18 TSMC_28 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_YDEC3TO8
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_YDEC3TO8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
XI32 TSMC_3 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI35 TSMC_6 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_3 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI38 TSMC_6 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI39 TSMC_3 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_19 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI42 TSMC_6 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI43 TSMC_3 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_6 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI33 VSS VSS TSMC_15 TSMC_13 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI34 VSS VSS TSMC_16 TSMC_12 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI37 VSS VSS TSMC_17 TSMC_11 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI40 VSS VSS TSMC_18 TSMC_10 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI41 VSS VSS TSMC_19 TSMC_9 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI44 VSS VSS TSMC_20 TSMC_8 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI29 VSS VSS TSMC_22 TSMC_14 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI45 VSS VSS TSMC_21 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WPREDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WPREDEC TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI VSS TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 
XXya TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 VDD VDDI VSS TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ S6ALLSVTFW40W20_RF_YDEC3TO8 
XXpb TSMC_5 TSMC_6 TSMC_13 TSMC_14 TSMC_27 TSMC_28 TSMC_29 TSMC_30 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DEC2TO4 
XXpd TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DEC2TO4 
XXpc TSMC_3 TSMC_4 TSMC_11 TSMC_12 TSMC_31 TSMC_32 TSMC_33 TSMC_34 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DEC2TO4 
XXpa TSMC_7 TSMC_8 TSMC_15 TSMC_16 TSMC_23 TSMC_24 TSMC_25 TSMC_26 VDD VDDI 
+ VSS S6ALLSVTFW40W20_RF_DECPDA 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ENLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_ENLAT TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS 
XI0 VSS VSS TSMC_1 TSMC_4 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI6 VSS VSS TSMC_5 TSMC_6 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI5 VSS VSS TSMC_4 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI4 VSS VSS TSMC_6 TSMC_3 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
MM5 TSMC_5 TSMC_6 TSMC_8 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_8 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_5 TSMC_2 TSMC_9 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_9 TSMC_4 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_5 TSMC_6 TSMC_10 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_10 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_5 TSMC_2 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_11 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WTUNE
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WTUNE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS TSMC_9 TSMC_10 TSMC_11 
XXenlat TSMC_1 TSMC_9 TSMC_8 VDD VDDI VSS S6ALLSVTFW40W20_RF_ENLAT 
XI15 VSS VSS TSMC_10 TSMC_11 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=7 n_l=0.020u p_totalM=3 p_nfin=7 p_l=0.020u 
XI9<2> VSS VSS TSMC_2 TSMC_12 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI9<1> VSS VSS TSMC_3 TSMC_13 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI9<0> VSS VSS TSMC_4 TSMC_14 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI8<2> VSS VSS TSMC_12 TSMC_5 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI8<1> VSS VSS TSMC_13 TSMC_6 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI8<0> VSS VSS TSMC_14 TSMC_7 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WPRCHBUF
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WPRCHBUF TSMC_1 TSMC_2 VDD VDDI VSS TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
XI18 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=7 p_l=0.020u 
XI17<7> TSMC_8 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<6> TSMC_9 TSMC_1 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<5> TSMC_10 TSMC_1 VSS VSS VDDI VDD TSMC_23 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<4> TSMC_11 TSMC_1 VSS VSS VDDI VDD TSMC_24 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<3> TSMC_4 TSMC_1 VSS VSS VDDI VDD TSMC_25 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<2> TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_26 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<1> TSMC_6 TSMC_1 VSS VSS VDDI VDD TSMC_27 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<0> TSMC_7 TSMC_1 VSS VSS VDDI VDD TSMC_28 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<7> TSMC_8 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<6> TSMC_9 TSMC_1 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<5> TSMC_10 TSMC_1 VSS VSS VDDI VDD TSMC_23 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<4> TSMC_11 TSMC_1 VSS VSS VDDI VDD TSMC_24 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<3> TSMC_4 TSMC_1 VSS VSS VDDI VDD TSMC_25 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<2> TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_26 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<1> TSMC_6 TSMC_1 VSS VSS VDDI VDD TSMC_27 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<0> TSMC_7 TSMC_1 VSS VSS VDDI VDD TSMC_28 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI7<7> VSS VSS TSMC_21 TSMC_12 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<6> VSS VSS TSMC_22 TSMC_13 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<5> VSS VSS TSMC_23 TSMC_14 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<4> VSS VSS TSMC_24 TSMC_15 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<3> VSS VSS TSMC_25 TSMC_16 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<2> VSS VSS TSMC_26 TSMC_17 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<1> VSS VSS TSMC_27 TSMC_18 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<0> VSS VSS TSMC_28 TSMC_19 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI2 VSS VSS TSMC_20 TSMC_3 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=9 n_l=16.0n p_totalM=6 p_nfin=9 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_ILATCH TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_svt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_svt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ADRLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_ADRLAT TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 VDD VDDI VSS 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 
XXylat<2> TSMC_33 TSMC_1 TSMC_2 TSMC_19 TSMC_22 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXylat<1> TSMC_34 TSMC_1 TSMC_2 TSMC_20 TSMC_23 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXylat<0> TSMC_35 TSMC_1 TSMC_2 TSMC_21 TSMC_24 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<7> TSMC_25 TSMC_1 TSMC_2 TSMC_3 TSMC_11 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<6> TSMC_26 TSMC_1 TSMC_2 TSMC_4 TSMC_12 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<5> TSMC_27 TSMC_1 TSMC_2 TSMC_5 TSMC_13 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<4> TSMC_28 TSMC_1 TSMC_2 TSMC_6 TSMC_14 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<3> TSMC_29 TSMC_1 TSMC_2 TSMC_7 TSMC_15 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<2> TSMC_30 TSMC_1 TSMC_2 TSMC_8 TSMC_16 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<1> TSMC_31 TSMC_1 TSMC_2 TSMC_9 TSMC_17 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
XXxlat<0> TSMC_32 TSMC_1 TSMC_2 TSMC_10 TSMC_18 VDD VDDI VSS 
+ S6ALLSVTFW40W20_ILATCH 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WGCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WGCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 VDD VDDI VSS TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 
XXclkgen TSMC_1 TSMC_33 TSMC_38 TSMC_62 TSMC_8 TSMC_9 TSMC_26 TSMC_31 VDD VDDI 
+ VSS TSMC_36 S6ALLSVTFW40W20_RF_WCLKGEN 
XXpredecs TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_10 TSMC_11 
+ TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 VDD VDDI VSS TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ S6ALLSVTFW40W20_RF_WPREDEC 
XXwtune TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_62 VDD VDDI VSS 
+ TSMC_32 TSMC_34 TSMC_35 S6ALLSVTFW40W20_RF_WTUNE 
XXwprchb TSMC_9 TSMC_26 VDD VDDI VSS TSMC_37 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 S6ALLSVTFW40W20_RF_WPRCHBUF 
XXadrlat TSMC_8 TSMC_9 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 VDD VDDI VSS 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 S6ALLSVTFW40W20_RF_ADRLAT 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_GCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_GCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 VDD VDDI VSS TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 
XXtiel TSMC_87 TSMC_88 VDD VSS S6ALLSVTFW40W20_RF_TIELGEN 
XXpudelay TSMC_27 TSMC_30 TSMC_86 VDD VSS S6ALLSVTFW40W20_RF_PUDELAY 
XXrctrl TSMC_1 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_20 
+ TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_29 TSMC_35 TSMC_36 TSMC_37 
+ TSMC_38 TSMC_71 TSMC_73 TSMC_89 TSMC_90 VDD VDDI VSS TSMC_75 TSMC_76 
+ TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 
+ TSMC_85 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 S6ALLSVTFW40W20_RF_RGCTRL 
XXdkctd TSMC_8 TSMC_9 TSMC_3 TSMC_13 TSMC_7 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_DKCTD 
XXwctrl TSMC_2 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_29 TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_89 VDD VDDI VSS 
+ TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 
+ S6ALLSVTFW40W20_RF_WGCTRL 
MM1_header VDDI TSMC_28 VDD VDD pch_svt_mac l=0.020u nfin=7 m=24 
XI13 VSS VSS TSMC_28 TSMC_139 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI29 VSS VSS TSMC_88 TSMC_140 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=6 n_l=0.020u p_totalM=1 
+ p_nfin=6 p_l=0.020u 
XI3 VSS VSS TSMC_140 TSMC_141 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=2 n_nfin=6 n_l=0.020u p_totalM=2 
+ p_nfin=6 p_l=0.020u 
XI12 VSS VSS TSMC_139 TSMC_29 VDD VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=8 n_nfin=5 n_l=0.020u p_totalM=8 
+ p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RCTD TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
XI79 TSMC_5 TSMC_6 VSS VSS VDDI VDD TSMC_7 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_2 TSMC_8 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_9 TSMC_6 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI76 TSMC_11 TSMC_10 VSS VSS VDDI VDD TSMC_4 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_12 TSMC_6 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI66 TSMC_2 TSMC_3 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_3 TSMC_15 VSS VSS VDDI VDD TSMC_5 
+ S6ALLSVTFW40W20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI149 VSS VSS TSMC_13 TSMC_16 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_11 TSMC_17 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI89 VSS VSS TSMC_14 TSMC_12 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_7 TSMC_18 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_19 TSMC_20 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_18 TSMC_8 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_21 TSMC_11 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_20 TSMC_15 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI145 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_11 TSMC_22 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI144 VSS VSS TSMC_23 TSMC_24 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI150 VSS VSS TSMC_13 TSMC_25 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_16 TSMC_23 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI143 VSS VSS TSMC_24 TSMC_19 VDDI VDD 
+ S6ALLSVTFW40W20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RDTRKEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_RDTRKEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS 
MM24 TSMC_11 TSMC_10 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM17 TSMC_4 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=4 m=4 
MM16 TSMC_4 TSMC_10 TSMC_12 VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM15 TSMC_12 TSMC_6 VSS VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM13 TSMC_3 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM8 TSMC_2 TSMC_10 TSMC_13 VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM2 TSMC_1 TSMC_14 TSMC_15 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM4 TSMC_15 TSMC_9 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM9 TSMC_16 TSMC_5 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM7 TSMC_13 TSMC_1 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM10 TSMC_3 TSMC_10 TSMC_16 VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM23 TSMC_2 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM3 VDDI TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM30 TSMC_10 TSMC_11 VDD VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM27 TSMC_2 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM20 TSMC_17 TSMC_6 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM19 TSMC_4 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=6 
MM18 TSMC_4 TSMC_11 TSMC_17 VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM14 TSMC_3 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM26 TSMC_3 TSMC_11 TSMC_18 VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM5 TSMC_19 TSMC_14 VDDI VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM0 TSMC_1 TSMC_14 TSMC_19 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM29 TSMC_2 TSMC_11 TSMC_20 VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM28 TSMC_20 TSMC_1 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM25 TSMC_18 TSMC_5 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM1 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.016u nfin=5 m=2 
XI33 TSMC_7 TSMC_2 TSMC_9 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW40W20_nand3_svt_mac_pcell n_totalM=2 n_nfin=6 n_l=0.016u p_totalM=2 
+ p_nfin=3 p_l=0.016u 
XI1 VSS VSS TSMC_1 TSMC_14 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKGIORD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TRKGIORD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 VDD VDDI VSS TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
XXrctd TSMC_4 TSMC_8 TSMC_9 TSMC_34 VDD VDDI VSS 
+ S6ALLSVTFW40W20_RF_RCTD 
XI23 VSS VSS TSMC_35 TSMC_36 VDDI VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI33 VSS VSS TSMC_18 TSMC_35 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XXrdtrken TSMC_4 TSMC_1 TSMC_2 TSMC_3 TSMC_5 TSMC_6 TSMC_34 TSMC_19 TSMC_36 
+ TSMC_20 TSMC_21 VDD VDDI VSS S6ALLSVTFW40W20_RF_RDTRKEN 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    16FF_2P_D130_v0d2_x1_for_BL_trk
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk TSMC_1 TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 VDD VSS TSMC_6 TSMC_7 TSMC_8 
MNpg_rp TSMC_3 TSMC_5 TSMC_9 VSS nchpg_8trpsr_mac l=20n nfin=2 m=1 
MNpd_rp TSMC_9 TSMC_1 VSS VSS nchpd_8trpsr_mac l=20n nfin=2 m=1 
MNpg_R TSMC_6 TSMC_8 TSMC_10 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MNpd_R TSMC_10 TSMC_11 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpd_L TSMC_11 TSMC_1 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpg_L TSMC_7 VSS TSMC_11 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MPpu_R TSMC_12 TSMC_11 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
MPpu_L TSMC_11 TSMC_1 TSMC_2 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    16FF_2P_D130_v0d2_x1_for_BL_trk_x2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 TSMC_1 TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 
XI1 TSMC_1 TSMC_3 TSMC_4 TSMC_5 TSMC_7 VDD VSS TSMC_10 TSMC_11 TSMC_12 
+ S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk 
XI0 TSMC_1 TSMC_2 TSMC_4 TSMC_6 TSMC_8 VDD VSS TSMC_9 TSMC_11 TSMC_13 
+ S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RBL_TRK_4X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_D130_ARRAY_RBL_TRK_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 VDD VDDAI 
+ VSS TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 
XI4 VDDAI TSMC_22 TSMC_5 TSMC_6 TSMC_8 TSMC_9 TSMC_12 TSMC_13 VDD VSS 
+ TSMC_23 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
+ S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
XI5 VDDAI TSMC_4 TSMC_22 TSMC_6 TSMC_10 TSMC_11 VSS VSS VDD VSS TSMC_15 
+ TSMC_23 TSMC_17 TSMC_20 TSMC_21 
+ S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WL_TRACK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_WL_TRACK TSMC_1 VSS TSMC_2 TSMC_3 
MMRWL VSS TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MMWWL1 VSS TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MMWWL0q VSS TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RWL_TRK_X2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 VDD VDDAI VSS TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
XI4 TSMC_5 VSS TSMC_5 TSMC_12 S6ALLSVTFW40W20_RF_WL_TRACK 
XI5 TSMC_5 VSS TSMC_5 TSMC_12 S6ALLSVTFW40W20_RF_WL_TRACK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PIN_GCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_PIN_GCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 VSS TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 
XD40 VSS TSMC_77 ndio_mac nfin=2 l=200.0n m=1 
XD39 VSS TSMC_49 ndio_mac nfin=2 l=200.0n m=1 
XD34 VSS TSMC_88 ndio_mac nfin=2 l=200.0n m=1 
XD41 VSS TSMC_78 ndio_mac nfin=2 l=200.0n m=1 
XD5<10> VSS TSMC_12 ndio_mac nfin=2 l=200.0n m=1 
XD5<9> VSS TSMC_13 ndio_mac nfin=2 l=200.0n m=1 
XD5<8> VSS TSMC_14 ndio_mac nfin=2 l=200.0n m=1 
XD5<7> VSS TSMC_15 ndio_mac nfin=2 l=200.0n m=1 
XD5<6> VSS TSMC_16 ndio_mac nfin=2 l=200.0n m=1 
XD5<5> VSS TSMC_17 ndio_mac nfin=2 l=200.0n m=1 
XD5<4> VSS TSMC_18 ndio_mac nfin=2 l=200.0n m=1 
XD5<3> VSS TSMC_19 ndio_mac nfin=2 l=200.0n m=1 
XD5<2> VSS TSMC_20 ndio_mac nfin=2 l=200.0n m=1 
XD5<1> VSS TSMC_21 ndio_mac nfin=2 l=200.0n m=1 
XD5<0> VSS TSMC_22 ndio_mac nfin=2 l=200.0n m=1 
XD8 VSS TSMC_81 ndio_mac nfin=2 l=200.0n m=1 
XD4<10> VSS TSMC_34 ndio_mac nfin=2 l=200.0n m=1 
XD4<9> VSS TSMC_35 ndio_mac nfin=2 l=200.0n m=1 
XD4<8> VSS TSMC_36 ndio_mac nfin=2 l=200.0n m=1 
XD4<7> VSS TSMC_37 ndio_mac nfin=2 l=200.0n m=1 
XD4<6> VSS TSMC_38 ndio_mac nfin=2 l=200.0n m=1 
XD4<5> VSS TSMC_39 ndio_mac nfin=2 l=200.0n m=1 
XD4<4> VSS TSMC_40 ndio_mac nfin=2 l=200.0n m=1 
XD4<3> VSS TSMC_41 ndio_mac nfin=2 l=200.0n m=1 
XD4<2> VSS TSMC_42 ndio_mac nfin=2 l=200.0n m=1 
XD4<1> VSS TSMC_43 ndio_mac nfin=2 l=200.0n m=1 
XD4<0> VSS TSMC_44 ndio_mac nfin=2 l=200.0n m=1 
XD25 VSS TSMC_48 ndio_mac nfin=2 l=200.0n m=1 
XD31<2> VSS TSMC_67 ndio_mac nfin=2 l=200.0n m=1 
XD31<1> VSS TSMC_68 ndio_mac nfin=2 l=200.0n m=1 
XD31<0> VSS TSMC_69 ndio_mac nfin=2 l=200.0n m=1 
XD21 VSS TSMC_92 ndio_mac nfin=2 l=200.0n m=1 
XD35<1> VSS TSMC_51 ndio_mac nfin=2 l=200.0n m=1 
XD35<0> VSS TSMC_52 ndio_mac nfin=2 l=200.0n m=1 
XDdummy<0> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<1> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<2> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<3> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<4> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<5> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD30<2> VSS TSMC_64 ndio_mac nfin=2 l=200.0n m=1 
XD30<1> VSS TSMC_65 ndio_mac nfin=2 l=200.0n m=1 
XD30<0> VSS TSMC_66 ndio_mac nfin=2 l=200.0n m=1 
XD28 VSS TSMC_47 ndio_mac nfin=2 l=200.0n m=1 
XD7 VSS TSMC_76 ndio_mac nfin=2 l=200.0n m=1 
XD2<10> VSS TSMC_23 ndio_mac nfin=2 l=200.0n m=1 
XD2<9> VSS TSMC_24 ndio_mac nfin=2 l=200.0n m=1 
XD2<8> VSS TSMC_25 ndio_mac nfin=2 l=200.0n m=1 
XD2<7> VSS TSMC_26 ndio_mac nfin=2 l=200.0n m=1 
XD2<6> VSS TSMC_27 ndio_mac nfin=2 l=200.0n m=1 
XD2<5> VSS TSMC_28 ndio_mac nfin=2 l=200.0n m=1 
XD2<4> VSS TSMC_29 ndio_mac nfin=2 l=200.0n m=1 
XD2<3> VSS TSMC_30 ndio_mac nfin=2 l=200.0n m=1 
XD2<2> VSS TSMC_31 ndio_mac nfin=2 l=200.0n m=1 
XD2<1> VSS TSMC_32 ndio_mac nfin=2 l=200.0n m=1 
XD2<0> VSS TSMC_33 ndio_mac nfin=2 l=200.0n m=1 
XD3<10> VSS TSMC_1 ndio_mac nfin=2 l=200.0n m=1 
XD3<9> VSS TSMC_2 ndio_mac nfin=2 l=200.0n m=1 
XD3<8> VSS TSMC_3 ndio_mac nfin=2 l=200.0n m=1 
XD3<7> VSS TSMC_4 ndio_mac nfin=2 l=200.0n m=1 
XD3<6> VSS TSMC_5 ndio_mac nfin=2 l=200.0n m=1 
XD3<5> VSS TSMC_6 ndio_mac nfin=2 l=200.0n m=1 
XD3<4> VSS TSMC_7 ndio_mac nfin=2 l=200.0n m=1 
XD3<3> VSS TSMC_8 ndio_mac nfin=2 l=200.0n m=1 
XD3<2> VSS TSMC_9 ndio_mac nfin=2 l=200.0n m=1 
XD3<1> VSS TSMC_10 ndio_mac nfin=2 l=200.0n m=1 
XD3<0> VSS TSMC_11 ndio_mac nfin=2 l=200.0n m=1 
XD0<1> VSS TSMC_71 ndio_mac nfin=2 l=200.0n m=1 
XD0<0> VSS TSMC_72 ndio_mac nfin=2 l=200.0n m=1 
XD24 VSS TSMC_46 ndio_mac nfin=2 l=200.0n m=1 
XD26 VSS TSMC_45 ndio_mac nfin=2 l=200.0n m=1 
XD6 VSS TSMC_50 ndio_mac nfin=2 l=200.0n m=1 
XD9 VSS TSMC_73 ndio_mac nfin=2 l=200.0n m=1 
XD20 VSS TSMC_91 ndio_mac nfin=2 l=200.0n m=1 
XD19 VSS TSMC_74 ndio_mac nfin=2 l=200.0n m=1 
XD38<8> VSS TSMC_53 ndio_mac nfin=2 l=200.0n m=1 
XD38<7> VSS TSMC_54 ndio_mac nfin=2 l=200.0n m=1 
XD38<6> VSS TSMC_55 ndio_mac nfin=2 l=200.0n m=1 
XD38<5> VSS TSMC_56 ndio_mac nfin=2 l=200.0n m=1 
XD38<4> VSS TSMC_57 ndio_mac nfin=2 l=200.0n m=1 
XD38<3> VSS TSMC_58 ndio_mac nfin=2 l=200.0n m=1 
XD38<2> VSS TSMC_59 ndio_mac nfin=2 l=200.0n m=1 
XD38<1> VSS TSMC_60 ndio_mac nfin=2 l=200.0n m=1 
XD38<0> VSS TSMC_61 ndio_mac nfin=2 l=200.0n m=1 
XD37 VSS TSMC_75 ndio_mac nfin=2 l=200.0n m=1 
XD42<1> VSS TSMC_79 ndio_mac nfin=2 l=200.0n m=1 
XD42<0> VSS TSMC_80 ndio_mac nfin=2 l=200.0n m=1 
XD1<1> VSS TSMC_89 ndio_mac nfin=2 l=200.0n m=1 
XD1<0> VSS TSMC_90 ndio_mac nfin=2 l=200.0n m=1 
XD29 VSS TSMC_87 ndio_mac nfin=2 l=200.0n m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    N16_2PRF_BITCELL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_N16_2PRF_BITCELL TSMC_1 TSMC_2 TSMC_3 VDD VSS TSMC_4 
+ TSMC_5 TSMC_6 
MNpg_rp TSMC_2 TSMC_3 TSMC_7 VSS nchpg_8trpsr_mac l=20n nfin=2 m=1 
MNpd_rp TSMC_7 TSMC_8 VSS VSS nchpd_8trpsr_mac l=20n nfin=2 m=1 
MNpd_L TSMC_9 TSMC_8 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpd_R TSMC_8 TSMC_9 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpg_R TSMC_5 TSMC_6 TSMC_8 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MNpg_L TSMC_4 TSMC_6 TSMC_9 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MPpu_L TSMC_9 TSMC_8 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
MPpu_R TSMC_8 TSMC_9 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_4X2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_D130_ARRAY_4X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 VDD VDDAI VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ TSMC_14 TSMC_15 TSMC_16 
XI7 VDDAI TSMC_3 TSMC_7 VDD VSS TSMC_9 TSMC_11 TSMC_15 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
XI6 VDDAI TSMC_4 TSMC_8 VDD VSS TSMC_10 TSMC_12 TSMC_16 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
XI5 VDDAI TSMC_3 TSMC_8 VDD VSS TSMC_9 TSMC_11 TSMC_16 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
XI4 VDDAI TSMC_4 TSMC_7 VDD VSS TSMC_10 TSMC_12 TSMC_15 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
XI3 VDDAI TSMC_4 TSMC_6 VDD VSS TSMC_10 TSMC_12 TSMC_14 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
XI2 VDDAI TSMC_3 TSMC_6 VDD VSS TSMC_9 TSMC_11 TSMC_14 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
XI1 VDDAI TSMC_4 TSMC_5 VDD VSS TSMC_10 TSMC_12 TSMC_13 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
XI0 VDDAI TSMC_3 TSMC_5 VDD VSS TSMC_9 TSMC_11 TSMC_13 
+ S6ALLSVTFW40W20_N16_2PRF_BITCELL 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RBL_TRK_OFF_4X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_D130_ARRAY_RBL_TRK_OFF_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDAI VSS TSMC_12 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
XI2 VDDAI TSMC_4 TSMC_20 TSMC_6 TSMC_10 TSMC_11 VSS VSS VDD VSS TSMC_12 
+ TSMC_21 TSMC_15 TSMC_18 TSMC_19 
+ S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
XI4 VDDAI TSMC_20 TSMC_5 TSMC_6 TSMC_8 TSMC_9 VSS VSS VDD VSS TSMC_21 
+ TSMC_13 TSMC_15 TSMC_16 TSMC_17 
+ S6ALLSVTFW40W20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RWL_TRK_X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X1 TSMC_1 TSMC_2 TSMC_3 VDD VDDAI 
+ VSS TSMC_4 TSMC_5 TSMC_6 TSMC_7 
XI2 TSMC_3 VSS TSMC_3 TSMC_7 S6ALLSVTFW40W20_RF_WL_TRACK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    LIO_PWR_TK_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_LIO_PWR_TK_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI 
+ TSMC_5 
MM_TKPKP3 TSMC_6 TSMC_3 TSMC_7 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP2 TSMC_7 TSMC_3 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP4 TSMC_5 TSMC_4 TSMC_6 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP1 TSMC_6 TSMC_2 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKLIO_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TRKLIO_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS 
MM0 TSMC_3 TSMC_4 VSS VSS nch_lvt_mac l=0.020u nfin=7 m=2 
MM5 TSMC_11 TSMC_9 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_1 TSMC_9 TSMC_11 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_9 TSMC_1 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM8 TSMC_12 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_9 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=2 
MM11 VDD TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_9 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=2 
MM7 TSMC_14 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM13 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM14 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_9 TSMC_1 TSMC_14 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI13 TSMC_5 TSMC_6 TSMC_7 TSMC_10 VDD VDDI TSMC_13 
+ S6ALLSVTFW40W20_LIO_PWR_TK_SVT_V1 
XXpwd0 TSMC_5 TSMC_6 TSMC_7 TSMC_10 VDD VDDI TSMC_13 
+ S6ALLSVTFW40W20_LIO_PWR_TK_SVT_V1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKLIOX2_72_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_TRKLIOX2_72_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 VDD VDDAI VDDI VSS TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 
XI35 VSS VSS TSMC_25 TSMC_26 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI31 VSS VSS TSMC_27 TSMC_28 VDD VDD S6ALLSVTFW40W20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XXtrklio TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_9 TSMC_10 TSMC_11 TSMC_26 TSMC_15 
+ TSMC_18 VDD VDDI VSS S6ALLSVTFW40W20_RF_TRKLIO_SVT_V1 
XI32 TSMC_14 TSMC_1 VSS VSS VDD VDD TSMC_27 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI38 TSMC_28 TSMC_16 VSS VSS VDD VDD TSMC_25 
+ S6ALLSVTFW40W20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    LIO_PWR_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_LIO_PWR_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI 
+ TSMC_5 
MM_PKP3 TSMC_5 TSMC_2 TSMC_6 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_PKP2 TSMC_6 TSMC_2 TSMC_7 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_PKP1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LIO_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_LIO_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 VDD VDDI VSS 
MM4 TSMC_1 TSMC_10 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM8 TSMC_11 TSMC_8 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_1 TSMC_7 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_2 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_2 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_13 TSMC_7 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI0 TSMC_4 TSMC_5 TSMC_6 TSMC_9 VDD VDD TSMC_12 
+ S6ALLSVTFW40W20_LIO_PWR_SVT_V1 
MM2 TSMC_3 TSMC_10 VSS VSS nch_lvt_mac l=0.020u nfin=7 m=2 
XI17 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW40W20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LIOX2_72_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_LIOX2_72_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDAI VDDI VSS 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 
XXlio0 TSMC_9 TSMC_11 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_12 
+ VDD VDDI VSS S6ALLSVTFW40W20_RF_LIO_SVT_V1 
XXlio1 TSMC_8 TSMC_10 TSMC_1 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_12 
+ VDD VDDI VSS S6ALLSVTFW40W20_RF_LIO_SVT_V1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PIN_GIO_MUX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VSS 
XD5 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD4 VSS TSMC_2 ndio_mac nfin=2 l=200.0n m=1 
XD6 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD1 VSS TSMC_3 ndio_mac nfin=2 l=200.0n m=1 
XD2 VSS TSMC_4 ndio_mac nfin=2 l=200.0n m=1 
XD3 VSS TSMC_1 ndio_mac nfin=2 l=200.0n m=1 
XD7 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<7> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<6> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<5> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<4> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<3> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<2> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<1> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD9<0> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD8 VSS VSS ndio_mac nfin=2 l=200.0n m=1 
.ENDS

.SUBCKT ndio_mac PLUS MINUS 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_inv_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_ulvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_inv_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_ulvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nand3_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_lvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nor2_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_ulvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nor2_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_lvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nand2_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_ulvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW40W20_nand2_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS





**** End of leaf cells

.SUBCKT S6ALLSVTFW40W20_PIN_ROW TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 VSS TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 
XPINIO0 TSMC_96 TSMC_210 TSMC_32 TSMC_178 TSMC_64 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO1 TSMC_95 TSMC_209 TSMC_31 TSMC_177 TSMC_63 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO2 TSMC_94 TSMC_208 TSMC_30 TSMC_176 TSMC_62 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO3 TSMC_93 TSMC_207 TSMC_29 TSMC_175 TSMC_61 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO4 TSMC_92 TSMC_206 TSMC_28 TSMC_174 TSMC_60 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO5 TSMC_91 TSMC_205 TSMC_27 TSMC_173 TSMC_59 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO6 TSMC_90 TSMC_204 TSMC_26 TSMC_172 TSMC_58 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO7 TSMC_89 TSMC_203 TSMC_25 TSMC_171 TSMC_57 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO8 TSMC_88 TSMC_202 TSMC_24 TSMC_170 TSMC_56 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO9 TSMC_87 TSMC_201 TSMC_23 TSMC_169 TSMC_55 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO10 TSMC_86 TSMC_200 TSMC_22 TSMC_168 TSMC_54 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO11 TSMC_85 TSMC_199 TSMC_21 TSMC_167 TSMC_53 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO12 TSMC_84 TSMC_198 TSMC_20 TSMC_166 TSMC_52 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO13 TSMC_83 TSMC_197 TSMC_19 TSMC_165 TSMC_51 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO14 TSMC_82 TSMC_196 TSMC_18 TSMC_164 TSMC_50 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO15 TSMC_81 TSMC_195 TSMC_17 TSMC_163 TSMC_49 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO16 TSMC_80 TSMC_194 TSMC_16 TSMC_162 TSMC_48 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO17 TSMC_79 TSMC_193 TSMC_15 TSMC_161 TSMC_47 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO18 TSMC_78 TSMC_192 TSMC_14 TSMC_160 TSMC_46 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO19 TSMC_77 TSMC_191 TSMC_13 TSMC_159 TSMC_45 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO20 TSMC_76 TSMC_190 TSMC_12 TSMC_158 TSMC_44 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO21 TSMC_75 TSMC_189 TSMC_11 TSMC_157 TSMC_43 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO22 TSMC_74 TSMC_188 TSMC_10 TSMC_156 TSMC_42 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO23 TSMC_73 TSMC_187 TSMC_9 TSMC_155 TSMC_41 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO24 TSMC_72 TSMC_186 TSMC_8 TSMC_154 TSMC_40 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO25 TSMC_71 TSMC_185 TSMC_7 TSMC_153 TSMC_39 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO26 TSMC_70 TSMC_184 TSMC_6 TSMC_152 TSMC_38 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO27 TSMC_69 TSMC_183 TSMC_5 TSMC_151 TSMC_37 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO28 TSMC_68 TSMC_182 TSMC_4 TSMC_150 TSMC_36 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO29 TSMC_67 TSMC_181 TSMC_3 TSMC_149 TSMC_35 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO30 TSMC_66 TSMC_180 TSMC_2 TSMC_148 TSMC_34 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINIO31 TSMC_65 TSMC_179 TSMC_1 TSMC_147 TSMC_33 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW40W20_RF_PIN_GIO_MUX4 
XPINCTRL TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_97 TSMC_98 TSMC_99 TSMC_100 
+ TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_136 
+ TSMC_235 TSMC_108 TSMC_121 TSMC_243 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 
+ TSMC_144 TSMC_145 TSMC_253 TSMC_254 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_236 TSMC_129 TSMC_130 TSMC_109 
+ TSMC_233 TSMC_146 TSMC_135 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_134 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_133 VSS TSMC_237 
+ TSMC_131 TSMC_132 TSMC_122 TSMC_234 S6ALLSVTFW40W20_RF_PIN_GCTRL 
.ENDS

.SUBCKT S6ALLSVTFW40W20_GCTRL_GIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 VDDI VDDM VSS TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 
+ TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 
+ TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 
+ TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 
+ TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 
+ TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 
+ TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 
+ TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 
+ TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 
+ TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 
+ TSMC_417 TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 
+ TSMC_425 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 
+ TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 
+ TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 
+ TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 
+ TSMC_473 TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 
+ TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 
+ TSMC_489 TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_504 
+ TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 
+ TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 
+ TSMC_521 TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 
+ TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 
+ TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 
+ TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 
+ TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 TSMC_567 TSMC_568 
+ TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 TSMC_578 TSMC_579 TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 
+ TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 
+ TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 TSMC_616 
+ TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 
+ TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 TSMC_631 TSMC_632 
+ TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 TSMC_639 TSMC_640 
+ TSMC_641 TSMC_642 TSMC_643 TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ TSMC_649 TSMC_650 TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 
+ TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 TSMC_664 
+ TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 TSMC_671 TSMC_672 
+ TSMC_673 TSMC_674 TSMC_675 TSMC_676 TSMC_677 TSMC_678 TSMC_679 TSMC_680 
+ TSMC_681 TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 TSMC_687 TSMC_688 
+ TSMC_689 TSMC_690 TSMC_691 TSMC_692 TSMC_693 TSMC_694 TSMC_695 TSMC_696 
+ TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_701 TSMC_702 TSMC_703 TSMC_704 
+ TSMC_705 TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 TSMC_711 TSMC_712 
+ TSMC_713 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 TSMC_719 TSMC_720 
+ TSMC_721 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_727 TSMC_728 
+ TSMC_729 TSMC_730 TSMC_731 TSMC_732 TSMC_733 TSMC_734 TSMC_735 TSMC_736 
+ TSMC_737 TSMC_738 TSMC_739 TSMC_740 TSMC_741 TSMC_742 TSMC_743 TSMC_744 
+ TSMC_745 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 TSMC_751 TSMC_752 
+ TSMC_753 TSMC_754 TSMC_755 TSMC_756 TSMC_757 TSMC_758 TSMC_759 TSMC_760 
+ TSMC_761 TSMC_762 TSMC_763 TSMC_764 TSMC_765 TSMC_766 TSMC_767 TSMC_768 
+ TSMC_769 TSMC_770 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_775 
XGIO_MUX0 TSMC_34 TSMC_66 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_742 TSMC_774 
+ TSMC_776 TSMC_242 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_646 TSMC_710 TSMC_678 TSMC_408 TSMC_409 
+ TSMC_410 TSMC_411 TSMC_536 TSMC_537 TSMC_538 TSMC_539 TSMC_574 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX1 TSMC_33 TSMC_65 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_741 TSMC_773 
+ TSMC_776 TSMC_241 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_645 TSMC_709 TSMC_677 TSMC_404 TSMC_405 
+ TSMC_406 TSMC_407 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_573 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX2 TSMC_32 TSMC_64 TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_740 TSMC_772 
+ TSMC_776 TSMC_240 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_644 TSMC_708 TSMC_676 TSMC_400 TSMC_401 
+ TSMC_402 TSMC_403 TSMC_528 TSMC_529 TSMC_530 TSMC_531 TSMC_572 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX3 TSMC_31 TSMC_63 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_739 TSMC_771 
+ TSMC_776 TSMC_239 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_643 TSMC_707 TSMC_675 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_571 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX4 TSMC_30 TSMC_62 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_738 TSMC_770 
+ TSMC_776 TSMC_238 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_642 TSMC_706 TSMC_674 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_570 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX5 TSMC_29 TSMC_61 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_737 TSMC_769 
+ TSMC_776 TSMC_237 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_641 TSMC_705 TSMC_673 TSMC_388 TSMC_389 
+ TSMC_390 TSMC_391 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_569 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX6 TSMC_28 TSMC_60 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_736 TSMC_768 
+ TSMC_776 TSMC_236 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_640 TSMC_704 TSMC_672 TSMC_384 TSMC_385 
+ TSMC_386 TSMC_387 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_568 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX7 TSMC_27 TSMC_59 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_735 TSMC_767 
+ TSMC_776 TSMC_235 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_639 TSMC_703 TSMC_671 TSMC_380 TSMC_381 
+ TSMC_382 TSMC_383 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_567 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX8 TSMC_26 TSMC_58 TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_734 TSMC_766 
+ TSMC_776 TSMC_234 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_638 TSMC_702 TSMC_670 TSMC_376 TSMC_377 
+ TSMC_378 TSMC_379 TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_566 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX9 TSMC_25 TSMC_57 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_733 TSMC_765 
+ TSMC_776 TSMC_233 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_637 TSMC_701 TSMC_669 TSMC_372 TSMC_373 
+ TSMC_374 TSMC_375 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_565 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX10 TSMC_24 TSMC_56 TSMC_151 TSMC_152 TSMC_153 TSMC_154 TSMC_732 
+ TSMC_764 TSMC_776 TSMC_232 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_636 TSMC_700 TSMC_668 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_496 TSMC_497 TSMC_498 TSMC_499 
+ TSMC_564 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX11 TSMC_23 TSMC_55 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_731 
+ TSMC_763 TSMC_776 TSMC_231 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_635 TSMC_699 TSMC_667 TSMC_364 
+ TSMC_365 TSMC_366 TSMC_367 TSMC_492 TSMC_493 TSMC_494 TSMC_495 
+ TSMC_563 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX12 TSMC_22 TSMC_54 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_730 
+ TSMC_762 TSMC_776 TSMC_230 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_634 TSMC_698 TSMC_666 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_488 TSMC_489 TSMC_490 TSMC_491 
+ TSMC_562 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX13 TSMC_21 TSMC_53 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_729 
+ TSMC_761 TSMC_776 TSMC_229 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_633 TSMC_697 TSMC_665 TSMC_356 
+ TSMC_357 TSMC_358 TSMC_359 TSMC_484 TSMC_485 TSMC_486 TSMC_487 
+ TSMC_561 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX14 TSMC_20 TSMC_52 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_728 
+ TSMC_760 TSMC_776 TSMC_228 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_632 TSMC_696 TSMC_664 TSMC_352 
+ TSMC_353 TSMC_354 TSMC_355 TSMC_480 TSMC_481 TSMC_482 TSMC_483 
+ TSMC_560 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX15 TSMC_19 TSMC_51 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_727 
+ TSMC_759 TSMC_776 TSMC_227 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_631 TSMC_695 TSMC_663 TSMC_348 
+ TSMC_349 TSMC_350 TSMC_351 TSMC_476 TSMC_477 TSMC_478 TSMC_479 
+ TSMC_559 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX16 TSMC_18 TSMC_50 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_726 
+ TSMC_758 TSMC_776 TSMC_226 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_630 TSMC_694 TSMC_662 TSMC_344 
+ TSMC_345 TSMC_346 TSMC_347 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_558 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX17 TSMC_17 TSMC_49 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_725 
+ TSMC_757 TSMC_776 TSMC_225 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_629 TSMC_693 TSMC_661 TSMC_340 
+ TSMC_341 TSMC_342 TSMC_343 TSMC_468 TSMC_469 TSMC_470 TSMC_471 
+ TSMC_557 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX18 TSMC_16 TSMC_48 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_724 
+ TSMC_756 TSMC_776 TSMC_224 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_628 TSMC_692 TSMC_660 TSMC_336 
+ TSMC_337 TSMC_338 TSMC_339 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_556 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX19 TSMC_15 TSMC_47 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_723 
+ TSMC_755 TSMC_776 TSMC_223 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_627 TSMC_691 TSMC_659 TSMC_332 
+ TSMC_333 TSMC_334 TSMC_335 TSMC_460 TSMC_461 TSMC_462 TSMC_463 
+ TSMC_555 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX20 TSMC_14 TSMC_46 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_722 
+ TSMC_754 TSMC_776 TSMC_222 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_626 TSMC_690 TSMC_658 TSMC_328 
+ TSMC_329 TSMC_330 TSMC_331 TSMC_456 TSMC_457 TSMC_458 TSMC_459 
+ TSMC_554 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX21 TSMC_13 TSMC_45 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_721 
+ TSMC_753 TSMC_776 TSMC_221 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_625 TSMC_689 TSMC_657 TSMC_324 
+ TSMC_325 TSMC_326 TSMC_327 TSMC_452 TSMC_453 TSMC_454 TSMC_455 
+ TSMC_553 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX22 TSMC_12 TSMC_44 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_720 
+ TSMC_752 TSMC_776 TSMC_220 TSMC_777 TSMC_778 TSMC_779 TSMC_780 
+ TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_624 TSMC_688 TSMC_656 TSMC_320 
+ TSMC_321 TSMC_322 TSMC_323 TSMC_448 TSMC_449 TSMC_450 TSMC_451 
+ TSMC_552 TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX23 TSMC_11 TSMC_43 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_719 
+ TSMC_751 TSMC_776 TSMC_219 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_623 TSMC_687 TSMC_655 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_551 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX24 TSMC_10 TSMC_42 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_718 
+ TSMC_750 TSMC_776 TSMC_218 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_622 TSMC_686 TSMC_654 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_550 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX25 TSMC_9 TSMC_41 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_717 
+ TSMC_749 TSMC_776 TSMC_217 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_621 TSMC_685 TSMC_653 TSMC_308 TSMC_309 
+ TSMC_310 TSMC_311 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_549 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX26 TSMC_8 TSMC_40 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_716 
+ TSMC_748 TSMC_776 TSMC_216 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_620 TSMC_684 TSMC_652 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_432 TSMC_433 TSMC_434 TSMC_435 TSMC_548 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX27 TSMC_7 TSMC_39 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_715 
+ TSMC_747 TSMC_776 TSMC_215 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_619 TSMC_683 TSMC_651 TSMC_300 TSMC_301 
+ TSMC_302 TSMC_303 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_547 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX28 TSMC_6 TSMC_38 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_714 
+ TSMC_746 TSMC_776 TSMC_214 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_618 TSMC_682 TSMC_650 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_424 TSMC_425 TSMC_426 TSMC_427 TSMC_546 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX29 TSMC_5 TSMC_37 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_713 
+ TSMC_745 TSMC_776 TSMC_213 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_617 TSMC_681 TSMC_649 TSMC_292 TSMC_293 
+ TSMC_294 TSMC_295 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_545 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX30 TSMC_4 TSMC_36 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_712 
+ TSMC_744 TSMC_776 TSMC_212 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_616 TSMC_680 TSMC_648 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_416 TSMC_417 TSMC_418 TSMC_419 TSMC_544 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XGIO_MUX31 TSMC_3 TSMC_35 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_711 
+ TSMC_743 TSMC_776 TSMC_211 TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 
+ TSMC_280 VDDM VDDI VSS TSMC_615 TSMC_679 TSMC_647 TSMC_284 TSMC_285 
+ TSMC_286 TSMC_287 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_543 
+ TSMC_782 TSMC_610 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_GIOM4 
XTRKGIOL TSMC_776 TSMC_787 TSMC_788 TSMC_789 TSMC_790 TSMC_777 TSMC_778 
+ TSMC_779 TSMC_780 TSMC_781 TSMC_280 VDDM VDDI VSS TSMC_791 TSMC_792 
+ TSMC_208 TSMC_540 TSMC_541 TSMC_209 TSMC_782 TSMC_610 TSMC_793 
+ TSMC_794 TSMC_795 TSMC_796 TSMC_797 TSMC_783 TSMC_784 TSMC_785 
+ TSMC_786 S6ALLSVTFW40W20_RF_TRKGIOWR 
XTRKGIOR TSMC_798 TSMC_798 TSMC_799 TSMC_195 TSMC_195 TSMC_281 TSMC_776 
+ TSMC_243 TSMC_244 TSMC_787 TSMC_788 TSMC_789 TSMC_790 TSMC_777 
+ TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_800 TSMC_281 TSMC_280 VDDM 
+ VDDI VSS TSMC_607 TSMC_801 TSMC_782 TSMC_610 TSMC_794 TSMC_795 
+ TSMC_796 TSMC_797 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ S6ALLSVTFW40W20_RF_TRKGIORD 
XGCTRL TSMC_1 TSMC_2 TSMC_612 TSMC_802 TSMC_613 TSMC_614 TSMC_611 TSMC_196 
+ TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_280 TSMC_803 TSMC_804 
+ TSMC_281 TSMC_805 TSMC_806 TSMC_807 TSMC_608 TSMC_210 TSMC_776 
+ TSMC_609 TSMC_808 TSMC_809 TSMC_810 TSMC_811 TSMC_245 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_812 TSMC_803 TSMC_804 TSMC_813 
+ TSMC_805 TSMC_806 TSMC_787 TSMC_788 TSMC_789 TSMC_790 TSMC_777 
+ TSMC_778 TSMC_779 TSMC_780 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 
+ TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_781 TSMC_267 TSMC_800 
+ TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 
+ TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_775 TSMC_281 
+ TSMC_280 TSMC_282 TSMC_283 VDDM VDDI VSS TSMC_542 TSMC_575 TSMC_576 TSMC_577 
+ TSMC_782 TSMC_578 TSMC_579 TSMC_580 TSMC_581 TSMC_582 TSMC_583 
+ TSMC_584 TSMC_585 TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 
+ TSMC_591 TSMC_592 TSMC_593 TSMC_594 TSMC_595 TSMC_610 TSMC_793 
+ TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 TSMC_602 
+ TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_794 TSMC_795 TSMC_796 TSMC_797 
+ TSMC_783 TSMC_784 TSMC_785 TSMC_786 TSMC_808 TSMC_809 TSMC_810 
+ TSMC_811 S6ALLSVTFW40W20_RF_GCTRL 
.ENDS

.SUBCKT S6ALLSVTFW40W20_ROW_TRACKING TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 
+ TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 
+ TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_377 
+ TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 VDDM 
+ VDDAI VDDI VSS TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 
XTRKROW0 TSMC_383 TSMC_384 TSMC_392 TSMC_393 TSMC_389 VDDM VDDAI VSS TSMC_127 
+ TSMC_128 TSMC_255 TSMC_256 TSMC_394 TSMC_395 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW1 TSMC_381 TSMC_382 TSMC_396 TSMC_397 TSMC_389 VDDM VDDAI VSS TSMC_125 
+ TSMC_126 TSMC_253 TSMC_254 TSMC_398 TSMC_399 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW2 TSMC_379 TSMC_380 TSMC_400 TSMC_401 TSMC_389 VDDM VDDAI VSS TSMC_123 
+ TSMC_124 TSMC_251 TSMC_252 TSMC_402 TSMC_403 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW3 TSMC_377 TSMC_378 TSMC_404 TSMC_405 TSMC_389 VDDM VDDAI VSS TSMC_121 
+ TSMC_122 TSMC_249 TSMC_250 TSMC_406 TSMC_407 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW4 TSMC_375 TSMC_376 TSMC_408 TSMC_409 TSMC_389 VDDM VDDAI VSS TSMC_119 
+ TSMC_120 TSMC_247 TSMC_248 TSMC_410 TSMC_411 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW5 TSMC_373 TSMC_374 TSMC_412 TSMC_413 TSMC_389 VDDM VDDAI VSS TSMC_117 
+ TSMC_118 TSMC_245 TSMC_246 TSMC_414 TSMC_415 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW6 TSMC_371 TSMC_372 TSMC_416 TSMC_417 TSMC_389 VDDM VDDAI VSS TSMC_115 
+ TSMC_116 TSMC_243 TSMC_244 TSMC_418 TSMC_419 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW7 TSMC_369 TSMC_370 TSMC_420 TSMC_421 TSMC_389 VDDM VDDAI VSS TSMC_113 
+ TSMC_114 TSMC_241 TSMC_242 TSMC_422 TSMC_423 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW8 TSMC_367 TSMC_368 TSMC_424 TSMC_425 TSMC_389 VDDM VDDAI VSS TSMC_111 
+ TSMC_112 TSMC_239 TSMC_240 TSMC_426 TSMC_427 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW9 TSMC_365 TSMC_366 TSMC_428 TSMC_429 TSMC_389 VDDM VDDAI VSS TSMC_109 
+ TSMC_110 TSMC_237 TSMC_238 TSMC_430 TSMC_431 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW10 TSMC_363 TSMC_364 TSMC_432 TSMC_433 TSMC_389 VDDM VDDAI VSS TSMC_107 
+ TSMC_108 TSMC_235 TSMC_236 TSMC_434 TSMC_435 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW11 TSMC_361 TSMC_362 TSMC_436 TSMC_437 TSMC_389 VDDM VDDAI VSS TSMC_105 
+ TSMC_106 TSMC_233 TSMC_234 TSMC_438 TSMC_439 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW12 TSMC_359 TSMC_360 TSMC_440 TSMC_441 TSMC_389 VDDM VDDAI VSS TSMC_103 
+ TSMC_104 TSMC_231 TSMC_232 TSMC_442 TSMC_443 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW13 TSMC_357 TSMC_358 TSMC_444 TSMC_445 TSMC_389 VDDM VDDAI VSS TSMC_101 
+ TSMC_102 TSMC_229 TSMC_230 TSMC_446 TSMC_447 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW14 TSMC_355 TSMC_356 TSMC_448 TSMC_449 TSMC_389 VDDM VDDAI VSS TSMC_99 
+ TSMC_100 TSMC_227 TSMC_228 TSMC_450 TSMC_451 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW15 TSMC_353 TSMC_354 TSMC_452 TSMC_453 TSMC_389 VDDM VDDAI VSS TSMC_97 
+ TSMC_98 TSMC_225 TSMC_226 TSMC_454 TSMC_455 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW16 TSMC_351 TSMC_352 TSMC_456 TSMC_457 TSMC_389 VDDM VDDAI VSS TSMC_95 
+ TSMC_96 TSMC_223 TSMC_224 TSMC_458 TSMC_459 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW17 TSMC_349 TSMC_350 TSMC_460 TSMC_461 TSMC_389 VDDM VDDAI VSS TSMC_93 
+ TSMC_94 TSMC_221 TSMC_222 TSMC_462 TSMC_463 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW18 TSMC_347 TSMC_348 TSMC_464 TSMC_465 TSMC_389 VDDM VDDAI VSS TSMC_91 
+ TSMC_92 TSMC_219 TSMC_220 TSMC_466 TSMC_467 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW19 TSMC_345 TSMC_346 TSMC_468 TSMC_469 TSMC_389 VDDM VDDAI VSS TSMC_89 
+ TSMC_90 TSMC_217 TSMC_218 TSMC_470 TSMC_471 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW20 TSMC_343 TSMC_344 TSMC_472 TSMC_473 TSMC_389 VDDM VDDAI VSS TSMC_87 
+ TSMC_88 TSMC_215 TSMC_216 TSMC_474 TSMC_475 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW21 TSMC_341 TSMC_342 TSMC_476 TSMC_477 TSMC_389 VDDM VDDAI VSS TSMC_85 
+ TSMC_86 TSMC_213 TSMC_214 TSMC_478 TSMC_479 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW22 TSMC_339 TSMC_340 TSMC_480 TSMC_481 TSMC_389 VDDM VDDAI VSS TSMC_83 
+ TSMC_84 TSMC_211 TSMC_212 TSMC_482 TSMC_483 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW23 TSMC_337 TSMC_338 TSMC_484 TSMC_485 TSMC_389 VDDM VDDAI VSS TSMC_81 
+ TSMC_82 TSMC_209 TSMC_210 TSMC_486 TSMC_487 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW24 TSMC_335 TSMC_336 TSMC_488 TSMC_489 TSMC_389 VDDM VDDAI VSS TSMC_79 
+ TSMC_80 TSMC_207 TSMC_208 TSMC_490 TSMC_491 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW25 TSMC_333 TSMC_334 TSMC_492 TSMC_493 TSMC_389 VDDM VDDAI VSS TSMC_77 
+ TSMC_78 TSMC_205 TSMC_206 TSMC_494 TSMC_495 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW26 TSMC_331 TSMC_332 TSMC_496 TSMC_497 TSMC_389 VDDM VDDAI VSS TSMC_75 
+ TSMC_76 TSMC_203 TSMC_204 TSMC_498 TSMC_499 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW27 TSMC_329 TSMC_330 TSMC_500 TSMC_501 TSMC_389 VDDM VDDAI VSS TSMC_73 
+ TSMC_74 TSMC_201 TSMC_202 TSMC_502 TSMC_503 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW28 TSMC_327 TSMC_328 TSMC_504 TSMC_505 TSMC_389 VDDM VDDAI VSS TSMC_71 
+ TSMC_72 TSMC_199 TSMC_200 TSMC_506 TSMC_507 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW29 TSMC_325 TSMC_326 TSMC_508 TSMC_509 TSMC_389 VDDM VDDAI VSS TSMC_69 
+ TSMC_70 TSMC_197 TSMC_198 TSMC_510 TSMC_511 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW30 TSMC_323 TSMC_324 TSMC_512 TSMC_513 TSMC_389 VDDM VDDAI VSS TSMC_67 
+ TSMC_68 TSMC_195 TSMC_196 TSMC_514 TSMC_515 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW31 TSMC_321 TSMC_322 TSMC_516 TSMC_517 TSMC_389 VDDM VDDAI VSS TSMC_65 
+ TSMC_66 TSMC_193 TSMC_194 TSMC_518 TSMC_519 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW32 TSMC_319 TSMC_320 TSMC_520 TSMC_521 TSMC_389 VDDM VDDAI VSS TSMC_63 
+ TSMC_64 TSMC_191 TSMC_192 TSMC_522 TSMC_523 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW33 TSMC_317 TSMC_318 TSMC_524 TSMC_525 TSMC_389 VDDM VDDAI VSS TSMC_61 
+ TSMC_62 TSMC_189 TSMC_190 TSMC_526 TSMC_527 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW34 TSMC_315 TSMC_316 TSMC_528 TSMC_529 TSMC_389 VDDM VDDAI VSS TSMC_59 
+ TSMC_60 TSMC_187 TSMC_188 TSMC_530 TSMC_531 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW35 TSMC_313 TSMC_314 TSMC_532 TSMC_533 TSMC_389 VDDM VDDAI VSS TSMC_57 
+ TSMC_58 TSMC_185 TSMC_186 TSMC_534 TSMC_535 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW36 TSMC_311 TSMC_312 TSMC_536 TSMC_537 TSMC_389 VDDM VDDAI VSS TSMC_55 
+ TSMC_56 TSMC_183 TSMC_184 TSMC_538 TSMC_539 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW37 TSMC_309 TSMC_310 TSMC_540 TSMC_541 TSMC_389 VDDM VDDAI VSS TSMC_53 
+ TSMC_54 TSMC_181 TSMC_182 TSMC_542 TSMC_543 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW38 TSMC_307 TSMC_308 TSMC_544 TSMC_545 TSMC_389 VDDM VDDAI VSS TSMC_51 
+ TSMC_52 TSMC_179 TSMC_180 TSMC_546 TSMC_547 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW39 TSMC_305 TSMC_306 TSMC_548 TSMC_549 TSMC_389 VDDM VDDAI VSS TSMC_49 
+ TSMC_50 TSMC_177 TSMC_178 TSMC_550 TSMC_551 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW40 TSMC_303 TSMC_304 TSMC_552 TSMC_553 TSMC_389 VDDM VDDAI VSS TSMC_47 
+ TSMC_48 TSMC_175 TSMC_176 TSMC_554 TSMC_555 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW41 TSMC_301 TSMC_302 TSMC_556 TSMC_557 TSMC_389 VDDM VDDAI VSS TSMC_45 
+ TSMC_46 TSMC_173 TSMC_174 TSMC_558 TSMC_559 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW42 TSMC_299 TSMC_300 TSMC_560 TSMC_561 TSMC_389 VDDM VDDAI VSS TSMC_43 
+ TSMC_44 TSMC_171 TSMC_172 TSMC_562 TSMC_563 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW43 TSMC_297 TSMC_298 TSMC_564 TSMC_565 TSMC_389 VDDM VDDAI VSS TSMC_41 
+ TSMC_42 TSMC_169 TSMC_170 TSMC_566 TSMC_567 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW44 TSMC_295 TSMC_296 TSMC_568 TSMC_569 TSMC_389 VDDM VDDAI VSS TSMC_39 
+ TSMC_40 TSMC_167 TSMC_168 TSMC_570 TSMC_571 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW45 TSMC_293 TSMC_294 TSMC_572 TSMC_573 TSMC_389 VDDM VDDAI VSS TSMC_37 
+ TSMC_38 TSMC_165 TSMC_166 TSMC_574 TSMC_575 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW46 TSMC_291 TSMC_292 TSMC_576 TSMC_577 TSMC_389 VDDM VDDAI VSS TSMC_35 
+ TSMC_36 TSMC_163 TSMC_164 TSMC_578 TSMC_579 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW47 TSMC_289 TSMC_290 TSMC_580 TSMC_581 TSMC_389 VDDM VDDAI VSS TSMC_33 
+ TSMC_34 TSMC_161 TSMC_162 TSMC_582 TSMC_583 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW48 TSMC_287 TSMC_288 TSMC_584 TSMC_585 TSMC_389 VDDM VDDAI VSS TSMC_31 
+ TSMC_32 TSMC_159 TSMC_160 TSMC_586 TSMC_587 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW49 TSMC_285 TSMC_286 TSMC_588 TSMC_589 TSMC_389 VDDM VDDAI VSS TSMC_29 
+ TSMC_30 TSMC_157 TSMC_158 TSMC_590 TSMC_591 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW50 TSMC_283 TSMC_284 TSMC_592 TSMC_593 TSMC_389 VDDM VDDAI VSS 
+ TSMC_27 TSMC_28 TSMC_155 TSMC_156 TSMC_594 TSMC_595 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW51 TSMC_281 TSMC_282 TSMC_596 TSMC_597 TSMC_389 VDDM VDDAI VSS 
+ TSMC_25 TSMC_26 TSMC_153 TSMC_154 TSMC_598 TSMC_599 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW52 TSMC_279 TSMC_280 TSMC_600 TSMC_601 TSMC_389 VDDM VDDAI VSS 
+ TSMC_23 TSMC_24 TSMC_151 TSMC_152 TSMC_602 TSMC_603 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW53 TSMC_277 TSMC_278 TSMC_604 TSMC_605 TSMC_389 VDDM VDDAI VSS 
+ TSMC_21 TSMC_22 TSMC_149 TSMC_150 TSMC_606 TSMC_607 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW54 TSMC_275 TSMC_276 TSMC_608 TSMC_609 TSMC_389 VDDM VDDAI VSS 
+ TSMC_19 TSMC_20 TSMC_147 TSMC_148 TSMC_610 TSMC_611 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW55 TSMC_273 TSMC_274 TSMC_612 TSMC_613 TSMC_389 VDDM VDDAI VSS 
+ TSMC_17 TSMC_18 TSMC_145 TSMC_146 TSMC_614 TSMC_615 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW56 TSMC_271 TSMC_272 TSMC_616 TSMC_617 TSMC_389 VDDM VDDAI VSS 
+ TSMC_15 TSMC_16 TSMC_143 TSMC_144 TSMC_618 TSMC_619 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW57 TSMC_269 TSMC_270 TSMC_620 TSMC_621 TSMC_389 VDDM VDDAI VSS 
+ TSMC_13 TSMC_14 TSMC_141 TSMC_142 TSMC_622 TSMC_623 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW58 TSMC_267 TSMC_268 TSMC_624 TSMC_625 TSMC_389 VDDM VDDAI VSS 
+ TSMC_11 TSMC_12 TSMC_139 TSMC_140 TSMC_626 TSMC_627 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW59 TSMC_265 TSMC_266 TSMC_628 TSMC_629 TSMC_389 VDDM VDDAI VSS 
+ TSMC_9 TSMC_10 TSMC_137 TSMC_138 TSMC_630 TSMC_631 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW60 TSMC_263 TSMC_264 TSMC_632 TSMC_633 TSMC_389 VDDM VDDAI VSS 
+ TSMC_7 TSMC_8 TSMC_135 TSMC_136 TSMC_634 TSMC_635 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW61 TSMC_261 TSMC_262 TSMC_636 TSMC_637 TSMC_389 VDDM VDDAI VSS 
+ TSMC_5 TSMC_6 TSMC_133 TSMC_134 TSMC_638 TSMC_639 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW62 TSMC_259 TSMC_260 TSMC_640 TSMC_641 TSMC_389 VDDM VDDAI VSS 
+ TSMC_3 TSMC_4 TSMC_131 TSMC_132 TSMC_642 TSMC_643 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROW63 TSMC_257 TSMC_258 TSMC_644 TSMC_645 TSMC_389 VDDM VDDAI VSS 
+ TSMC_1 TSMC_2 TSMC_129 TSMC_130 TSMC_646 TSMC_647 VSS 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XTRKROWL TSMC_648 TSMC_649 TSMC_389 VDDM VDDAI VSS TSMC_390 TSMC_650 
+ TSMC_651 VSS S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X1 
XTRKROWR TSMC_385 TSMC_652 TSMC_389 VDDM VDDAI VSS TSMC_391 TSMC_653 
+ TSMC_654 VSS S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X1 
XTRKCTRL TSMC_655 TSMC_656 TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 
+ TSMC_662 TSMC_663 TSMC_664 TSMC_665 TSMC_388 TSMC_386 TSMC_387 
+ TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 TSMC_671 TSMC_672 
+ TSMC_673 TSMC_674 TSMC_675 TSMC_676 TSMC_677 TSMC_678 TSMC_679 
+ TSMC_680 TSMC_681 TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 TSMC_687 
+ TSMC_389 VDDM VDDI VSS TSMC_688 TSMC_689 TSMC_690 TSMC_691 TSMC_692 
+ TSMC_693 TSMC_694 TSMC_695 TSMC_696 TSMC_697 TSMC_698 TSMC_699 
+ TSMC_700 TSMC_701 TSMC_702 TSMC_703 TSMC_704 TSMC_705 
+ S6ALLSVTFW40W20_RF_TRKCTRL 
.ENDS

.SUBCKT S6ALLSVTFW40W20_ARY4ROW TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 
+ TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 
+ TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_377 
+ TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 
+ TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 
+ TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 
+ TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 
+ TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 
+ TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_441 
+ TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_449 
+ TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_457 
+ TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 
+ TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 
+ TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 
+ TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_497 
+ TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_505 
+ TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_513 
+ TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_521 
+ TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 
+ TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 VDDM VDDAI 
+ VDDI VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 
+ TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 
+ TSMC_552 TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 TSMC_567 
XCOL0 TSMC_127 TSMC_128 TSMC_255 TSMC_256 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_383 TSMC_384 TSMC_511 TSMC_512 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL1 TSMC_125 TSMC_126 TSMC_253 TSMC_254 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_381 TSMC_382 TSMC_509 TSMC_510 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL2 TSMC_123 TSMC_124 TSMC_251 TSMC_252 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_379 TSMC_380 TSMC_507 TSMC_508 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL3 TSMC_121 TSMC_122 TSMC_249 TSMC_250 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_377 TSMC_378 TSMC_505 TSMC_506 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL4 TSMC_119 TSMC_120 TSMC_247 TSMC_248 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_375 TSMC_376 TSMC_503 TSMC_504 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL5 TSMC_117 TSMC_118 TSMC_245 TSMC_246 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_373 TSMC_374 TSMC_501 TSMC_502 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL6 TSMC_115 TSMC_116 TSMC_243 TSMC_244 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_371 TSMC_372 TSMC_499 TSMC_500 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL7 TSMC_113 TSMC_114 TSMC_241 TSMC_242 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_369 TSMC_370 TSMC_497 TSMC_498 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL8 TSMC_111 TSMC_112 TSMC_239 TSMC_240 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_367 TSMC_368 TSMC_495 TSMC_496 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL9 TSMC_109 TSMC_110 TSMC_237 TSMC_238 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_365 TSMC_366 TSMC_493 TSMC_494 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL10 TSMC_107 TSMC_108 TSMC_235 TSMC_236 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_363 TSMC_364 TSMC_491 TSMC_492 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL11 TSMC_105 TSMC_106 TSMC_233 TSMC_234 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_361 TSMC_362 TSMC_489 TSMC_490 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL12 TSMC_103 TSMC_104 TSMC_231 TSMC_232 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_359 TSMC_360 TSMC_487 TSMC_488 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL13 TSMC_101 TSMC_102 TSMC_229 TSMC_230 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_357 TSMC_358 TSMC_485 TSMC_486 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL14 TSMC_99 TSMC_100 TSMC_227 TSMC_228 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_355 TSMC_356 TSMC_483 TSMC_484 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL15 TSMC_97 TSMC_98 TSMC_225 TSMC_226 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_353 TSMC_354 TSMC_481 TSMC_482 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL16 TSMC_95 TSMC_96 TSMC_223 TSMC_224 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_351 TSMC_352 TSMC_479 TSMC_480 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL17 TSMC_93 TSMC_94 TSMC_221 TSMC_222 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_349 TSMC_350 TSMC_477 TSMC_478 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL18 TSMC_91 TSMC_92 TSMC_219 TSMC_220 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_347 TSMC_348 TSMC_475 TSMC_476 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL19 TSMC_89 TSMC_90 TSMC_217 TSMC_218 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_345 TSMC_346 TSMC_473 TSMC_474 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL20 TSMC_87 TSMC_88 TSMC_215 TSMC_216 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_343 TSMC_344 TSMC_471 TSMC_472 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL21 TSMC_85 TSMC_86 TSMC_213 TSMC_214 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_341 TSMC_342 TSMC_469 TSMC_470 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL22 TSMC_83 TSMC_84 TSMC_211 TSMC_212 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_339 TSMC_340 TSMC_467 TSMC_468 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL23 TSMC_81 TSMC_82 TSMC_209 TSMC_210 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_337 TSMC_338 TSMC_465 TSMC_466 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL24 TSMC_79 TSMC_80 TSMC_207 TSMC_208 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_335 TSMC_336 TSMC_463 TSMC_464 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL25 TSMC_77 TSMC_78 TSMC_205 TSMC_206 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_333 TSMC_334 TSMC_461 TSMC_462 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL26 TSMC_75 TSMC_76 TSMC_203 TSMC_204 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_331 TSMC_332 TSMC_459 TSMC_460 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL27 TSMC_73 TSMC_74 TSMC_201 TSMC_202 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_329 TSMC_330 TSMC_457 TSMC_458 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL28 TSMC_71 TSMC_72 TSMC_199 TSMC_200 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_327 TSMC_328 TSMC_455 TSMC_456 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL29 TSMC_69 TSMC_70 TSMC_197 TSMC_198 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_325 TSMC_326 TSMC_453 TSMC_454 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL30 TSMC_67 TSMC_68 TSMC_195 TSMC_196 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_323 TSMC_324 TSMC_451 TSMC_452 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL31 TSMC_65 TSMC_66 TSMC_193 TSMC_194 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_321 TSMC_322 TSMC_449 TSMC_450 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL32 TSMC_63 TSMC_64 TSMC_191 TSMC_192 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_319 TSMC_320 TSMC_447 TSMC_448 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL33 TSMC_61 TSMC_62 TSMC_189 TSMC_190 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_317 TSMC_318 TSMC_445 TSMC_446 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL34 TSMC_59 TSMC_60 TSMC_187 TSMC_188 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_315 TSMC_316 TSMC_443 TSMC_444 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL35 TSMC_57 TSMC_58 TSMC_185 TSMC_186 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_313 TSMC_314 TSMC_441 TSMC_442 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL36 TSMC_55 TSMC_56 TSMC_183 TSMC_184 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_311 TSMC_312 TSMC_439 TSMC_440 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL37 TSMC_53 TSMC_54 TSMC_181 TSMC_182 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_309 TSMC_310 TSMC_437 TSMC_438 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL38 TSMC_51 TSMC_52 TSMC_179 TSMC_180 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_307 TSMC_308 TSMC_435 TSMC_436 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL39 TSMC_49 TSMC_50 TSMC_177 TSMC_178 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_305 TSMC_306 TSMC_433 TSMC_434 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL40 TSMC_47 TSMC_48 TSMC_175 TSMC_176 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_303 TSMC_304 TSMC_431 TSMC_432 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL41 TSMC_45 TSMC_46 TSMC_173 TSMC_174 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_301 TSMC_302 TSMC_429 TSMC_430 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL42 TSMC_43 TSMC_44 TSMC_171 TSMC_172 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_299 TSMC_300 TSMC_427 TSMC_428 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL43 TSMC_41 TSMC_42 TSMC_169 TSMC_170 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_297 TSMC_298 TSMC_425 TSMC_426 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL44 TSMC_39 TSMC_40 TSMC_167 TSMC_168 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_295 TSMC_296 TSMC_423 TSMC_424 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL45 TSMC_37 TSMC_38 TSMC_165 TSMC_166 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_293 TSMC_294 TSMC_421 TSMC_422 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL46 TSMC_35 TSMC_36 TSMC_163 TSMC_164 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_291 TSMC_292 TSMC_419 TSMC_420 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL47 TSMC_33 TSMC_34 TSMC_161 TSMC_162 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_289 TSMC_290 TSMC_417 TSMC_418 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL48 TSMC_31 TSMC_32 TSMC_159 TSMC_160 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_287 TSMC_288 TSMC_415 TSMC_416 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL49 TSMC_29 TSMC_30 TSMC_157 TSMC_158 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_285 TSMC_286 TSMC_413 TSMC_414 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL50 TSMC_27 TSMC_28 TSMC_155 TSMC_156 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_283 TSMC_284 TSMC_411 TSMC_412 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL51 TSMC_25 TSMC_26 TSMC_153 TSMC_154 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_281 TSMC_282 TSMC_409 TSMC_410 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL52 TSMC_23 TSMC_24 TSMC_151 TSMC_152 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_279 TSMC_280 TSMC_407 TSMC_408 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL53 TSMC_21 TSMC_22 TSMC_149 TSMC_150 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_277 TSMC_278 TSMC_405 TSMC_406 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL54 TSMC_19 TSMC_20 TSMC_147 TSMC_148 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_275 TSMC_276 TSMC_403 TSMC_404 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL55 TSMC_17 TSMC_18 TSMC_145 TSMC_146 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_273 TSMC_274 TSMC_401 TSMC_402 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL56 TSMC_15 TSMC_16 TSMC_143 TSMC_144 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_271 TSMC_272 TSMC_399 TSMC_400 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL57 TSMC_13 TSMC_14 TSMC_141 TSMC_142 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_269 TSMC_270 TSMC_397 TSMC_398 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL58 TSMC_11 TSMC_12 TSMC_139 TSMC_140 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_267 TSMC_268 TSMC_395 TSMC_396 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL59 TSMC_9 TSMC_10 TSMC_137 TSMC_138 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_265 TSMC_266 TSMC_393 TSMC_394 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL60 TSMC_7 TSMC_8 TSMC_135 TSMC_136 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_263 TSMC_264 TSMC_391 TSMC_392 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL61 TSMC_5 TSMC_6 TSMC_133 TSMC_134 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_261 TSMC_262 TSMC_389 TSMC_390 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL62 TSMC_3 TSMC_4 TSMC_131 TSMC_132 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_259 TSMC_260 TSMC_387 TSMC_388 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL63 TSMC_1 TSMC_2 TSMC_129 TSMC_130 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ VDDM VDDAI VSS TSMC_257 TSMC_258 TSMC_385 TSMC_386 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XTRKL TSMC_513 TSMC_576 TSMC_577 TSMC_564 TSMC_565 TSMC_514 TSMC_514 
+ TSMC_568 TSMC_569 TSMC_570 TSMC_571 VDDM VDDAI VSS TSMC_560 TSMC_561 VSS 
+ TSMC_515 TSMC_572 TSMC_573 TSMC_574 TSMC_575 
+ S6ALLSVTFW40W20_D130_ARRAY_RBL_TRK_OFF_4X1 
XTRKR TSMC_516 TSMC_578 TSMC_579 TSMC_566 TSMC_567 TSMC_514 TSMC_514 
+ TSMC_568 TSMC_569 TSMC_570 TSMC_571 VDDM VDDAI VSS TSMC_562 TSMC_563 VSS 
+ TSMC_517 TSMC_572 TSMC_573 TSMC_574 TSMC_575 
+ S6ALLSVTFW40W20_D130_ARRAY_RBL_TRK_OFF_4X1 
XDEC TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_518 TSMC_518 TSMC_519 TSMC_520 TSMC_521 
+ TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 
+ TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_568 
+ TSMC_569 TSMC_570 TSMC_571 TSMC_536 VDDM VDDI VDDI VSS TSMC_537 
+ TSMC_538 TSMC_539 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 
+ TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 
+ TSMC_551 TSMC_552 TSMC_553 TSMC_554 TSMC_555 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ S6ALLSVTFW40W20_RF_XDEC4 
.ENDS

.SUBCKT S6ALLSVTFW40W20_ARY4ROW_TK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 
+ TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 
+ TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_377 
+ TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 
+ TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 
+ TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 
+ TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 
+ TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 
+ TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_441 
+ TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_449 
+ TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_457 
+ TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 
+ TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 
+ TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 
+ TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_497 
+ TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_505 
+ TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_513 
+ TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_521 
+ TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 
+ TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 VDDM VDDAI 
+ VDDI VSS TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 
+ TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 
+ TSMC_552 TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 TSMC_567 
+ TSMC_568 TSMC_569 
XCOL0 TSMC_127 TSMC_128 TSMC_255 TSMC_256 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_383 TSMC_384 TSMC_511 TSMC_512 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL1 TSMC_125 TSMC_126 TSMC_253 TSMC_254 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_381 TSMC_382 TSMC_509 TSMC_510 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL2 TSMC_123 TSMC_124 TSMC_251 TSMC_252 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_379 TSMC_380 TSMC_507 TSMC_508 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL3 TSMC_121 TSMC_122 TSMC_249 TSMC_250 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_377 TSMC_378 TSMC_505 TSMC_506 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL4 TSMC_119 TSMC_120 TSMC_247 TSMC_248 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_375 TSMC_376 TSMC_503 TSMC_504 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL5 TSMC_117 TSMC_118 TSMC_245 TSMC_246 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_373 TSMC_374 TSMC_501 TSMC_502 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL6 TSMC_115 TSMC_116 TSMC_243 TSMC_244 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_371 TSMC_372 TSMC_499 TSMC_500 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL7 TSMC_113 TSMC_114 TSMC_241 TSMC_242 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_369 TSMC_370 TSMC_497 TSMC_498 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL8 TSMC_111 TSMC_112 TSMC_239 TSMC_240 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_367 TSMC_368 TSMC_495 TSMC_496 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL9 TSMC_109 TSMC_110 TSMC_237 TSMC_238 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_365 TSMC_366 TSMC_493 TSMC_494 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL10 TSMC_107 TSMC_108 TSMC_235 TSMC_236 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_363 TSMC_364 TSMC_491 TSMC_492 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL11 TSMC_105 TSMC_106 TSMC_233 TSMC_234 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_361 TSMC_362 TSMC_489 TSMC_490 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL12 TSMC_103 TSMC_104 TSMC_231 TSMC_232 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_359 TSMC_360 TSMC_487 TSMC_488 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL13 TSMC_101 TSMC_102 TSMC_229 TSMC_230 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_357 TSMC_358 TSMC_485 TSMC_486 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL14 TSMC_99 TSMC_100 TSMC_227 TSMC_228 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_355 TSMC_356 TSMC_483 TSMC_484 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL15 TSMC_97 TSMC_98 TSMC_225 TSMC_226 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_353 TSMC_354 TSMC_481 TSMC_482 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL16 TSMC_95 TSMC_96 TSMC_223 TSMC_224 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_351 TSMC_352 TSMC_479 TSMC_480 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL17 TSMC_93 TSMC_94 TSMC_221 TSMC_222 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_349 TSMC_350 TSMC_477 TSMC_478 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL18 TSMC_91 TSMC_92 TSMC_219 TSMC_220 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_347 TSMC_348 TSMC_475 TSMC_476 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL19 TSMC_89 TSMC_90 TSMC_217 TSMC_218 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_345 TSMC_346 TSMC_473 TSMC_474 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL20 TSMC_87 TSMC_88 TSMC_215 TSMC_216 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_343 TSMC_344 TSMC_471 TSMC_472 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL21 TSMC_85 TSMC_86 TSMC_213 TSMC_214 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_341 TSMC_342 TSMC_469 TSMC_470 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL22 TSMC_83 TSMC_84 TSMC_211 TSMC_212 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_339 TSMC_340 TSMC_467 TSMC_468 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL23 TSMC_81 TSMC_82 TSMC_209 TSMC_210 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_337 TSMC_338 TSMC_465 TSMC_466 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL24 TSMC_79 TSMC_80 TSMC_207 TSMC_208 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_335 TSMC_336 TSMC_463 TSMC_464 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL25 TSMC_77 TSMC_78 TSMC_205 TSMC_206 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_333 TSMC_334 TSMC_461 TSMC_462 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL26 TSMC_75 TSMC_76 TSMC_203 TSMC_204 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_331 TSMC_332 TSMC_459 TSMC_460 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL27 TSMC_73 TSMC_74 TSMC_201 TSMC_202 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_329 TSMC_330 TSMC_457 TSMC_458 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL28 TSMC_71 TSMC_72 TSMC_199 TSMC_200 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_327 TSMC_328 TSMC_455 TSMC_456 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL29 TSMC_69 TSMC_70 TSMC_197 TSMC_198 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_325 TSMC_326 TSMC_453 TSMC_454 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL30 TSMC_67 TSMC_68 TSMC_195 TSMC_196 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_323 TSMC_324 TSMC_451 TSMC_452 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL31 TSMC_65 TSMC_66 TSMC_193 TSMC_194 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_321 TSMC_322 TSMC_449 TSMC_450 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL32 TSMC_63 TSMC_64 TSMC_191 TSMC_192 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_319 TSMC_320 TSMC_447 TSMC_448 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL33 TSMC_61 TSMC_62 TSMC_189 TSMC_190 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_317 TSMC_318 TSMC_445 TSMC_446 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL34 TSMC_59 TSMC_60 TSMC_187 TSMC_188 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_315 TSMC_316 TSMC_443 TSMC_444 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL35 TSMC_57 TSMC_58 TSMC_185 TSMC_186 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_313 TSMC_314 TSMC_441 TSMC_442 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL36 TSMC_55 TSMC_56 TSMC_183 TSMC_184 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_311 TSMC_312 TSMC_439 TSMC_440 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL37 TSMC_53 TSMC_54 TSMC_181 TSMC_182 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_309 TSMC_310 TSMC_437 TSMC_438 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL38 TSMC_51 TSMC_52 TSMC_179 TSMC_180 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_307 TSMC_308 TSMC_435 TSMC_436 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL39 TSMC_49 TSMC_50 TSMC_177 TSMC_178 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_305 TSMC_306 TSMC_433 TSMC_434 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL40 TSMC_47 TSMC_48 TSMC_175 TSMC_176 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_303 TSMC_304 TSMC_431 TSMC_432 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL41 TSMC_45 TSMC_46 TSMC_173 TSMC_174 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_301 TSMC_302 TSMC_429 TSMC_430 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL42 TSMC_43 TSMC_44 TSMC_171 TSMC_172 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_299 TSMC_300 TSMC_427 TSMC_428 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL43 TSMC_41 TSMC_42 TSMC_169 TSMC_170 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_297 TSMC_298 TSMC_425 TSMC_426 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL44 TSMC_39 TSMC_40 TSMC_167 TSMC_168 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_295 TSMC_296 TSMC_423 TSMC_424 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL45 TSMC_37 TSMC_38 TSMC_165 TSMC_166 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_293 TSMC_294 TSMC_421 TSMC_422 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL46 TSMC_35 TSMC_36 TSMC_163 TSMC_164 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_291 TSMC_292 TSMC_419 TSMC_420 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL47 TSMC_33 TSMC_34 TSMC_161 TSMC_162 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_289 TSMC_290 TSMC_417 TSMC_418 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL48 TSMC_31 TSMC_32 TSMC_159 TSMC_160 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_287 TSMC_288 TSMC_415 TSMC_416 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL49 TSMC_29 TSMC_30 TSMC_157 TSMC_158 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_285 TSMC_286 TSMC_413 TSMC_414 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL50 TSMC_27 TSMC_28 TSMC_155 TSMC_156 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_283 TSMC_284 TSMC_411 TSMC_412 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL51 TSMC_25 TSMC_26 TSMC_153 TSMC_154 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_281 TSMC_282 TSMC_409 TSMC_410 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL52 TSMC_23 TSMC_24 TSMC_151 TSMC_152 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_279 TSMC_280 TSMC_407 TSMC_408 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL53 TSMC_21 TSMC_22 TSMC_149 TSMC_150 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_277 TSMC_278 TSMC_405 TSMC_406 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL54 TSMC_19 TSMC_20 TSMC_147 TSMC_148 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_275 TSMC_276 TSMC_403 TSMC_404 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL55 TSMC_17 TSMC_18 TSMC_145 TSMC_146 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_273 TSMC_274 TSMC_401 TSMC_402 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL56 TSMC_15 TSMC_16 TSMC_143 TSMC_144 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_271 TSMC_272 TSMC_399 TSMC_400 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL57 TSMC_13 TSMC_14 TSMC_141 TSMC_142 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_269 TSMC_270 TSMC_397 TSMC_398 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL58 TSMC_11 TSMC_12 TSMC_139 TSMC_140 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_267 TSMC_268 TSMC_395 TSMC_396 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL59 TSMC_9 TSMC_10 TSMC_137 TSMC_138 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_265 TSMC_266 TSMC_393 TSMC_394 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL60 TSMC_7 TSMC_8 TSMC_135 TSMC_136 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_263 TSMC_264 TSMC_391 TSMC_392 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL61 TSMC_5 TSMC_6 TSMC_133 TSMC_134 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_261 TSMC_262 TSMC_389 TSMC_390 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL62 TSMC_3 TSMC_4 TSMC_131 TSMC_132 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_259 TSMC_260 TSMC_387 TSMC_388 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XCOL63 TSMC_1 TSMC_2 TSMC_129 TSMC_130 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ VDDM VDDAI VSS TSMC_257 TSMC_258 TSMC_385 TSMC_386 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_4X2 
XTRKL TSMC_513 TSMC_578 TSMC_579 TSMC_566 TSMC_567 TSMC_514 TSMC_514 
+ TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_564 TSMC_564 VDDM VDDAI VSS VSS 
+ TSMC_560 TSMC_561 TSMC_515 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_RBL_TRK_4X1 
XTRKR TSMC_580 TSMC_581 TSMC_582 TSMC_568 TSMC_569 TSMC_514 TSMC_514 
+ TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_565 TSMC_565 VDDM VDDAI VSS VSS 
+ TSMC_562 TSMC_563 TSMC_517 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 S6ALLSVTFW40W20_D130_ARRAY_RBL_TRK_4X1 
XDEC TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 
+ TSMC_591 TSMC_592 TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 
+ TSMC_598 TSMC_599 TSMC_518 TSMC_518 TSMC_519 TSMC_520 TSMC_521 
+ TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 
+ TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_570 
+ TSMC_571 TSMC_572 TSMC_573 TSMC_536 VDDM VDDI VDDI VSS TSMC_537 
+ TSMC_538 TSMC_539 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 
+ TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 
+ TSMC_551 TSMC_552 TSMC_553 TSMC_554 TSMC_555 TSMC_574 TSMC_575 TSMC_576 
+ TSMC_577 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ S6ALLSVTFW40W20_RF_XDEC4 
.ENDS

.SUBCKT S6ALLSVTFW40W20_LIO_LCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 
+ TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 
+ TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_377 
+ TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 
+ TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 
+ TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 
+ TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 
+ TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 
+ TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_441 
+ TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_449 
+ TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_457 
+ TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 
+ TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 
+ TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 
+ TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_497 
+ TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_505 
+ TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_513 
+ TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_521 
+ TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 
+ TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 
+ TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 
+ TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 TSMC_561 
+ TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 TSMC_567 TSMC_568 TSMC_569 
+ TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 TSMC_575 TSMC_576 TSMC_577 
+ TSMC_578 TSMC_579 TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 
+ TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 
+ TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 TSMC_609 
+ TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 
+ TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 TSMC_625 
+ TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 TSMC_631 TSMC_632 TSMC_633 
+ TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 
+ TSMC_642 TSMC_643 TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 
+ TSMC_650 TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 TSMC_657 
+ TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 TSMC_664 TSMC_665 
+ TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 TSMC_671 TSMC_672 TSMC_673 
+ TSMC_674 TSMC_675 TSMC_676 TSMC_677 TSMC_678 TSMC_679 TSMC_680 TSMC_681 
+ TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 TSMC_687 TSMC_688 TSMC_689 
+ TSMC_690 TSMC_691 TSMC_692 TSMC_693 TSMC_694 TSMC_695 VDDM VDDI VDDAI VSS 
+ TSMC_696 TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_701 TSMC_702 TSMC_703 
+ TSMC_704 TSMC_705 TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 TSMC_711 
+ TSMC_712 TSMC_713 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 TSMC_719 
+ TSMC_720 TSMC_721 
XLIO0 TSMC_127 TSMC_128 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_255 
+ TSMC_256 TSMC_383 TSMC_384 TSMC_693 VDDM VDDAI VDDI VSS TSMC_511 
+ TSMC_512 TSMC_639 TSMC_640 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO1 TSMC_125 TSMC_126 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_253 
+ TSMC_254 TSMC_381 TSMC_382 TSMC_693 VDDM VDDAI VDDI VSS TSMC_509 
+ TSMC_510 TSMC_637 TSMC_638 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO2 TSMC_123 TSMC_124 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_251 
+ TSMC_252 TSMC_379 TSMC_380 TSMC_693 VDDM VDDAI VDDI VSS TSMC_507 
+ TSMC_508 TSMC_635 TSMC_636 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO3 TSMC_121 TSMC_122 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_249 
+ TSMC_250 TSMC_377 TSMC_378 TSMC_693 VDDM VDDAI VDDI VSS TSMC_505 
+ TSMC_506 TSMC_633 TSMC_634 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO4 TSMC_119 TSMC_120 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_247 
+ TSMC_248 TSMC_375 TSMC_376 TSMC_693 VDDM VDDAI VDDI VSS TSMC_503 
+ TSMC_504 TSMC_631 TSMC_632 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO5 TSMC_117 TSMC_118 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_245 
+ TSMC_246 TSMC_373 TSMC_374 TSMC_693 VDDM VDDAI VDDI VSS TSMC_501 
+ TSMC_502 TSMC_629 TSMC_630 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO6 TSMC_115 TSMC_116 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_243 
+ TSMC_244 TSMC_371 TSMC_372 TSMC_693 VDDM VDDAI VDDI VSS TSMC_499 
+ TSMC_500 TSMC_627 TSMC_628 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO7 TSMC_113 TSMC_114 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_241 
+ TSMC_242 TSMC_369 TSMC_370 TSMC_693 VDDM VDDAI VDDI VSS TSMC_497 
+ TSMC_498 TSMC_625 TSMC_626 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO8 TSMC_111 TSMC_112 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_239 
+ TSMC_240 TSMC_367 TSMC_368 TSMC_693 VDDM VDDAI VDDI VSS TSMC_495 
+ TSMC_496 TSMC_623 TSMC_624 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO9 TSMC_109 TSMC_110 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 TSMC_237 
+ TSMC_238 TSMC_365 TSMC_366 TSMC_693 VDDM VDDAI VDDI VSS TSMC_493 
+ TSMC_494 TSMC_621 TSMC_622 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO10 TSMC_107 TSMC_108 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_235 TSMC_236 TSMC_363 TSMC_364 TSMC_693 VDDM VDDAI VDDI VSS TSMC_491 
+ TSMC_492 TSMC_619 TSMC_620 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO11 TSMC_105 TSMC_106 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_233 TSMC_234 TSMC_361 TSMC_362 TSMC_693 VDDM VDDAI VDDI VSS TSMC_489 
+ TSMC_490 TSMC_617 TSMC_618 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO12 TSMC_103 TSMC_104 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_231 TSMC_232 TSMC_359 TSMC_360 TSMC_693 VDDM VDDAI VDDI VSS TSMC_487 
+ TSMC_488 TSMC_615 TSMC_616 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO13 TSMC_101 TSMC_102 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_229 TSMC_230 TSMC_357 TSMC_358 TSMC_693 VDDM VDDAI VDDI VSS TSMC_485 
+ TSMC_486 TSMC_613 TSMC_614 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO14 TSMC_99 TSMC_100 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_227 TSMC_228 TSMC_355 TSMC_356 TSMC_693 VDDM VDDAI VDDI VSS TSMC_483 
+ TSMC_484 TSMC_611 TSMC_612 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO15 TSMC_97 TSMC_98 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_225 TSMC_226 TSMC_353 TSMC_354 TSMC_693 VDDM VDDAI VDDI VSS TSMC_481 
+ TSMC_482 TSMC_609 TSMC_610 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO16 TSMC_95 TSMC_96 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_223 TSMC_224 TSMC_351 TSMC_352 TSMC_693 VDDM VDDAI VDDI VSS TSMC_479 
+ TSMC_480 TSMC_607 TSMC_608 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO17 TSMC_93 TSMC_94 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_221 TSMC_222 TSMC_349 TSMC_350 TSMC_693 VDDM VDDAI VDDI VSS TSMC_477 
+ TSMC_478 TSMC_605 TSMC_606 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO18 TSMC_91 TSMC_92 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_219 TSMC_220 TSMC_347 TSMC_348 TSMC_693 VDDM VDDAI VDDI VSS TSMC_475 
+ TSMC_476 TSMC_603 TSMC_604 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO19 TSMC_89 TSMC_90 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_217 TSMC_218 TSMC_345 TSMC_346 TSMC_693 VDDM VDDAI VDDI VSS TSMC_473 
+ TSMC_474 TSMC_601 TSMC_602 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO20 TSMC_87 TSMC_88 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_215 TSMC_216 TSMC_343 TSMC_344 TSMC_693 VDDM VDDAI VDDI VSS TSMC_471 
+ TSMC_472 TSMC_599 TSMC_600 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO21 TSMC_85 TSMC_86 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_213 TSMC_214 TSMC_341 TSMC_342 TSMC_693 VDDM VDDAI VDDI VSS TSMC_469 
+ TSMC_470 TSMC_597 TSMC_598 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO22 TSMC_83 TSMC_84 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_211 TSMC_212 TSMC_339 TSMC_340 TSMC_693 VDDM VDDAI VDDI VSS TSMC_467 
+ TSMC_468 TSMC_595 TSMC_596 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO23 TSMC_81 TSMC_82 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_209 TSMC_210 TSMC_337 TSMC_338 TSMC_693 VDDM VDDAI VDDI VSS TSMC_465 
+ TSMC_466 TSMC_593 TSMC_594 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO24 TSMC_79 TSMC_80 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_207 TSMC_208 TSMC_335 TSMC_336 TSMC_693 VDDM VDDAI VDDI VSS TSMC_463 
+ TSMC_464 TSMC_591 TSMC_592 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO25 TSMC_77 TSMC_78 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_205 TSMC_206 TSMC_333 TSMC_334 TSMC_693 VDDM VDDAI VDDI VSS TSMC_461 
+ TSMC_462 TSMC_589 TSMC_590 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO26 TSMC_75 TSMC_76 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_203 TSMC_204 TSMC_331 TSMC_332 TSMC_693 VDDM VDDAI VDDI VSS TSMC_459 
+ TSMC_460 TSMC_587 TSMC_588 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO27 TSMC_73 TSMC_74 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_201 TSMC_202 TSMC_329 TSMC_330 TSMC_693 VDDM VDDAI VDDI VSS TSMC_457 
+ TSMC_458 TSMC_585 TSMC_586 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO28 TSMC_71 TSMC_72 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_199 TSMC_200 TSMC_327 TSMC_328 TSMC_693 VDDM VDDAI VDDI VSS TSMC_455 
+ TSMC_456 TSMC_583 TSMC_584 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO29 TSMC_69 TSMC_70 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_197 TSMC_198 TSMC_325 TSMC_326 TSMC_693 VDDM VDDAI VDDI VSS TSMC_453 
+ TSMC_454 TSMC_581 TSMC_582 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO30 TSMC_67 TSMC_68 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_195 TSMC_196 TSMC_323 TSMC_324 TSMC_693 VDDM VDDAI VDDI VSS TSMC_451 
+ TSMC_452 TSMC_579 TSMC_580 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO31 TSMC_65 TSMC_66 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_193 TSMC_194 TSMC_321 TSMC_322 TSMC_693 VDDM VDDAI VDDI VSS TSMC_449 
+ TSMC_450 TSMC_577 TSMC_578 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO32 TSMC_63 TSMC_64 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_191 TSMC_192 TSMC_319 TSMC_320 TSMC_693 VDDM VDDAI VDDI VSS TSMC_447 
+ TSMC_448 TSMC_575 TSMC_576 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO33 TSMC_61 TSMC_62 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_189 TSMC_190 TSMC_317 TSMC_318 TSMC_693 VDDM VDDAI VDDI VSS TSMC_445 
+ TSMC_446 TSMC_573 TSMC_574 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO34 TSMC_59 TSMC_60 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_187 TSMC_188 TSMC_315 TSMC_316 TSMC_693 VDDM VDDAI VDDI VSS TSMC_443 
+ TSMC_444 TSMC_571 TSMC_572 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO35 TSMC_57 TSMC_58 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_185 TSMC_186 TSMC_313 TSMC_314 TSMC_693 VDDM VDDAI VDDI VSS TSMC_441 
+ TSMC_442 TSMC_569 TSMC_570 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO36 TSMC_55 TSMC_56 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_183 TSMC_184 TSMC_311 TSMC_312 TSMC_693 VDDM VDDAI VDDI VSS TSMC_439 
+ TSMC_440 TSMC_567 TSMC_568 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO37 TSMC_53 TSMC_54 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_181 TSMC_182 TSMC_309 TSMC_310 TSMC_693 VDDM VDDAI VDDI VSS TSMC_437 
+ TSMC_438 TSMC_565 TSMC_566 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO38 TSMC_51 TSMC_52 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_179 TSMC_180 TSMC_307 TSMC_308 TSMC_693 VDDM VDDAI VDDI VSS TSMC_435 
+ TSMC_436 TSMC_563 TSMC_564 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO39 TSMC_49 TSMC_50 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_177 TSMC_178 TSMC_305 TSMC_306 TSMC_693 VDDM VDDAI VDDI VSS TSMC_433 
+ TSMC_434 TSMC_561 TSMC_562 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO40 TSMC_47 TSMC_48 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_175 TSMC_176 TSMC_303 TSMC_304 TSMC_693 VDDM VDDAI VDDI VSS TSMC_431 
+ TSMC_432 TSMC_559 TSMC_560 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO41 TSMC_45 TSMC_46 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_173 TSMC_174 TSMC_301 TSMC_302 TSMC_693 VDDM VDDAI VDDI VSS TSMC_429 
+ TSMC_430 TSMC_557 TSMC_558 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO42 TSMC_43 TSMC_44 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_171 TSMC_172 TSMC_299 TSMC_300 TSMC_693 VDDM VDDAI VDDI VSS TSMC_427 
+ TSMC_428 TSMC_555 TSMC_556 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO43 TSMC_41 TSMC_42 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_169 TSMC_170 TSMC_297 TSMC_298 TSMC_693 VDDM VDDAI VDDI VSS TSMC_425 
+ TSMC_426 TSMC_553 TSMC_554 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO44 TSMC_39 TSMC_40 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_167 TSMC_168 TSMC_295 TSMC_296 TSMC_693 VDDM VDDAI VDDI VSS TSMC_423 
+ TSMC_424 TSMC_551 TSMC_552 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO45 TSMC_37 TSMC_38 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_165 TSMC_166 TSMC_293 TSMC_294 TSMC_693 VDDM VDDAI VDDI VSS TSMC_421 
+ TSMC_422 TSMC_549 TSMC_550 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO46 TSMC_35 TSMC_36 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_163 TSMC_164 TSMC_291 TSMC_292 TSMC_693 VDDM VDDAI VDDI VSS TSMC_419 
+ TSMC_420 TSMC_547 TSMC_548 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO47 TSMC_33 TSMC_34 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_161 TSMC_162 TSMC_289 TSMC_290 TSMC_693 VDDM VDDAI VDDI VSS TSMC_417 
+ TSMC_418 TSMC_545 TSMC_546 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO48 TSMC_31 TSMC_32 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_159 TSMC_160 TSMC_287 TSMC_288 TSMC_693 VDDM VDDAI VDDI VSS TSMC_415 
+ TSMC_416 TSMC_543 TSMC_544 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO49 TSMC_29 TSMC_30 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_157 TSMC_158 TSMC_285 TSMC_286 TSMC_693 VDDM VDDAI VDDI VSS TSMC_413 
+ TSMC_414 TSMC_541 TSMC_542 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO50 TSMC_27 TSMC_28 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_155 TSMC_156 TSMC_283 TSMC_284 TSMC_693 VDDM VDDAI VDDI VSS TSMC_411 
+ TSMC_412 TSMC_539 TSMC_540 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO51 TSMC_25 TSMC_26 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_153 TSMC_154 TSMC_281 TSMC_282 TSMC_693 VDDM VDDAI VDDI VSS TSMC_409 
+ TSMC_410 TSMC_537 TSMC_538 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO52 TSMC_23 TSMC_24 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_151 TSMC_152 TSMC_279 TSMC_280 TSMC_693 VDDM VDDAI VDDI VSS TSMC_407 
+ TSMC_408 TSMC_535 TSMC_536 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO53 TSMC_21 TSMC_22 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_149 TSMC_150 TSMC_277 TSMC_278 TSMC_693 VDDM VDDAI VDDI VSS TSMC_405 
+ TSMC_406 TSMC_533 TSMC_534 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO54 TSMC_19 TSMC_20 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_147 TSMC_148 TSMC_275 TSMC_276 TSMC_693 VDDM VDDAI VDDI VSS TSMC_403 
+ TSMC_404 TSMC_531 TSMC_532 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO55 TSMC_17 TSMC_18 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_145 TSMC_146 TSMC_273 TSMC_274 TSMC_693 VDDM VDDAI VDDI VSS TSMC_401 
+ TSMC_402 TSMC_529 TSMC_530 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO56 TSMC_15 TSMC_16 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_143 TSMC_144 TSMC_271 TSMC_272 TSMC_693 VDDM VDDAI VDDI VSS TSMC_399 
+ TSMC_400 TSMC_527 TSMC_528 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO57 TSMC_13 TSMC_14 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_141 TSMC_142 TSMC_269 TSMC_270 TSMC_693 VDDM VDDAI VDDI VSS TSMC_397 
+ TSMC_398 TSMC_525 TSMC_526 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO58 TSMC_11 TSMC_12 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_139 TSMC_140 TSMC_267 TSMC_268 TSMC_693 VDDM VDDAI VDDI VSS TSMC_395 
+ TSMC_396 TSMC_523 TSMC_524 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO59 TSMC_9 TSMC_10 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_137 TSMC_138 TSMC_265 TSMC_266 TSMC_693 VDDM VDDAI VDDI VSS TSMC_393 
+ TSMC_394 TSMC_521 TSMC_522 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO60 TSMC_7 TSMC_8 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_135 TSMC_136 TSMC_263 TSMC_264 TSMC_693 VDDM VDDAI VDDI VSS TSMC_391 
+ TSMC_392 TSMC_519 TSMC_520 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO61 TSMC_5 TSMC_6 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_133 TSMC_134 TSMC_261 TSMC_262 TSMC_693 VDDM VDDAI VDDI VSS TSMC_389 
+ TSMC_390 TSMC_517 TSMC_518 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO62 TSMC_3 TSMC_4 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_131 TSMC_132 TSMC_259 TSMC_260 TSMC_693 VDDM VDDAI VDDI VSS TSMC_387 
+ TSMC_388 TSMC_515 TSMC_516 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XLIO63 TSMC_1 TSMC_2 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_129 TSMC_130 TSMC_257 TSMC_258 TSMC_693 VDDM VDDAI VDDI VSS TSMC_385 
+ TSMC_386 TSMC_513 TSMC_514 S6ALLSVTFW40W20_RF_LIOX2_72_V1 
XTROLIOL TSMC_719 TSMC_641 TSMC_717 TSMC_642 TSMC_643 TSMC_722 TSMC_723 
+ TSMC_724 TSMC_727 TSMC_728 TSMC_729 TSMC_725 TSMC_726 TSMC_644 
+ TSMC_645 TSMC_721 TSMC_647 TSMC_693 VDDM VDDAI VDDI VSS TSMC_730 
+ TSMC_649 TSMC_731 TSMC_651 TSMC_652 TSMC_653 
+ S6ALLSVTFW40W20_RF_TRKLIOX2_72_V1 
XTROLIOR TSMC_719 TSMC_654 TSMC_732 TSMC_655 TSMC_656 TSMC_722 TSMC_723 
+ TSMC_724 TSMC_727 TSMC_728 TSMC_729 TSMC_725 TSMC_726 TSMC_644 
+ TSMC_645 TSMC_721 TSMC_657 TSMC_693 VDDM VDDAI VDDI VSS TSMC_658 
+ TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 
+ S6ALLSVTFW40W20_RF_TRKLIOX2_72_V1 
XLCTRL TSMC_718 TSMC_664 TSMC_665 TSMC_719 TSMC_720 TSMC_733 TSMC_734 TSMC_722 
+ TSMC_723 TSMC_724 TSMC_727 TSMC_728 TSMC_729 TSMC_666 TSMC_667 
+ TSMC_668 TSMC_669 TSMC_670 TSMC_671 TSMC_725 TSMC_726 TSMC_644 
+ TSMC_735 TSMC_672 TSMC_646 TSMC_673 TSMC_674 TSMC_675 TSMC_676 
+ TSMC_677 TSMC_678 TSMC_679 TSMC_680 TSMC_681 TSMC_682 TSMC_683 TSMC_684 
+ TSMC_685 TSMC_686 TSMC_687 TSMC_688 TSMC_689 TSMC_690 TSMC_691 
+ TSMC_692 TSMC_693 TSMC_645 TSMC_694 TSMC_695 VDDM VDDI VSS TSMC_696 
+ TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_701 TSMC_702 TSMC_703 
+ TSMC_704 TSMC_705 TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 
+ TSMC_711 TSMC_712 TSMC_713 TSMC_714 TSMC_715 TSMC_716 
+ S6ALLSVTFW40W20_RF_LCTRL 
.ENDS

.SUBCKT S6ALLSVTFW40W20_WRITE_TRAKING TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 
+ TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 
+ TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_377 
+ TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 
+ TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 
+ TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 
+ TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 
+ TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 
+ TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 
+ TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_441 
+ TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_449 
+ TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_457 
+ TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 
+ TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 
+ TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 
+ TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_497 
+ TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_505 
+ TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_513 
+ TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_521 
+ TSMC_522 TSMC_523 VDDM VDDI VDDAI VSS TSMC_524 TSMC_525 TSMC_526 TSMC_527 
+ TSMC_528 
XRWLLD0 TSMC_127 TSMC_128 TSMC_255 TSMC_256 VSS VDDM VDDAI VSS TSMC_511 
+ TSMC_512 TSMC_383 TSMC_384 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD1 TSMC_125 TSMC_126 TSMC_253 TSMC_254 VSS VDDM VDDAI VSS TSMC_509 
+ TSMC_510 TSMC_381 TSMC_382 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD2 TSMC_123 TSMC_124 TSMC_251 TSMC_252 VSS VDDM VDDAI VSS TSMC_507 
+ TSMC_508 TSMC_379 TSMC_380 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD3 TSMC_121 TSMC_122 TSMC_249 TSMC_250 VSS VDDM VDDAI VSS TSMC_505 
+ TSMC_506 TSMC_377 TSMC_378 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD4 TSMC_119 TSMC_120 TSMC_247 TSMC_248 VSS VDDM VDDAI VSS TSMC_503 
+ TSMC_504 TSMC_375 TSMC_376 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD5 TSMC_117 TSMC_118 TSMC_245 TSMC_246 VSS VDDM VDDAI VSS TSMC_501 
+ TSMC_502 TSMC_373 TSMC_374 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD6 TSMC_115 TSMC_116 TSMC_243 TSMC_244 VSS VDDM VDDAI VSS TSMC_499 
+ TSMC_500 TSMC_371 TSMC_372 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD7 TSMC_113 TSMC_114 TSMC_241 TSMC_242 VSS VDDM VDDAI VSS TSMC_497 
+ TSMC_498 TSMC_369 TSMC_370 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD8 TSMC_111 TSMC_112 TSMC_239 TSMC_240 VSS VDDM VDDAI VSS TSMC_495 
+ TSMC_496 TSMC_367 TSMC_368 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD9 TSMC_109 TSMC_110 TSMC_237 TSMC_238 VSS VDDM VDDAI VSS TSMC_493 
+ TSMC_494 TSMC_365 TSMC_366 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD10 TSMC_107 TSMC_108 TSMC_235 TSMC_236 VSS VDDM VDDAI VSS TSMC_491 
+ TSMC_492 TSMC_363 TSMC_364 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD11 TSMC_105 TSMC_106 TSMC_233 TSMC_234 VSS VDDM VDDAI VSS TSMC_489 
+ TSMC_490 TSMC_361 TSMC_362 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD12 TSMC_103 TSMC_104 TSMC_231 TSMC_232 VSS VDDM VDDAI VSS TSMC_487 
+ TSMC_488 TSMC_359 TSMC_360 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD13 TSMC_101 TSMC_102 TSMC_229 TSMC_230 VSS VDDM VDDAI VSS TSMC_485 
+ TSMC_486 TSMC_357 TSMC_358 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD14 TSMC_99 TSMC_100 TSMC_227 TSMC_228 VSS VDDM VDDAI VSS TSMC_483 
+ TSMC_484 TSMC_355 TSMC_356 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD15 TSMC_97 TSMC_98 TSMC_225 TSMC_226 VSS VDDM VDDAI VSS TSMC_481 
+ TSMC_482 TSMC_353 TSMC_354 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD16 TSMC_95 TSMC_96 TSMC_223 TSMC_224 VSS VDDM VDDAI VSS TSMC_479 
+ TSMC_480 TSMC_351 TSMC_352 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD17 TSMC_93 TSMC_94 TSMC_221 TSMC_222 VSS VDDM VDDAI VSS TSMC_477 
+ TSMC_478 TSMC_349 TSMC_350 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD18 TSMC_91 TSMC_92 TSMC_219 TSMC_220 VSS VDDM VDDAI VSS TSMC_475 
+ TSMC_476 TSMC_347 TSMC_348 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD19 TSMC_89 TSMC_90 TSMC_217 TSMC_218 VSS VDDM VDDAI VSS TSMC_473 
+ TSMC_474 TSMC_345 TSMC_346 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD20 TSMC_87 TSMC_88 TSMC_215 TSMC_216 VSS VDDM VDDAI VSS TSMC_471 
+ TSMC_472 TSMC_343 TSMC_344 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD21 TSMC_85 TSMC_86 TSMC_213 TSMC_214 VSS VDDM VDDAI VSS TSMC_469 
+ TSMC_470 TSMC_341 TSMC_342 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD22 TSMC_83 TSMC_84 TSMC_211 TSMC_212 VSS VDDM VDDAI VSS TSMC_467 
+ TSMC_468 TSMC_339 TSMC_340 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD23 TSMC_81 TSMC_82 TSMC_209 TSMC_210 VSS VDDM VDDAI VSS TSMC_465 
+ TSMC_466 TSMC_337 TSMC_338 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD24 TSMC_79 TSMC_80 TSMC_207 TSMC_208 VSS VDDM VDDAI VSS TSMC_463 
+ TSMC_464 TSMC_335 TSMC_336 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD25 TSMC_77 TSMC_78 TSMC_205 TSMC_206 VSS VDDM VDDAI VSS TSMC_461 
+ TSMC_462 TSMC_333 TSMC_334 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD26 TSMC_75 TSMC_76 TSMC_203 TSMC_204 VSS VDDM VDDAI VSS TSMC_459 
+ TSMC_460 TSMC_331 TSMC_332 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD27 TSMC_73 TSMC_74 TSMC_201 TSMC_202 VSS VDDM VDDAI VSS TSMC_457 
+ TSMC_458 TSMC_329 TSMC_330 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD28 TSMC_71 TSMC_72 TSMC_199 TSMC_200 VSS VDDM VDDAI VSS TSMC_455 
+ TSMC_456 TSMC_327 TSMC_328 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD29 TSMC_69 TSMC_70 TSMC_197 TSMC_198 VSS VDDM VDDAI VSS TSMC_453 
+ TSMC_454 TSMC_325 TSMC_326 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD30 TSMC_67 TSMC_68 TSMC_195 TSMC_196 VSS VDDM VDDAI VSS TSMC_451 
+ TSMC_452 TSMC_323 TSMC_324 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD31 TSMC_65 TSMC_66 TSMC_193 TSMC_194 VSS VDDM VDDAI VSS TSMC_449 
+ TSMC_450 TSMC_321 TSMC_322 TSMC_529 TSMC_530 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD32 TSMC_63 TSMC_64 TSMC_191 TSMC_192 VSS VDDM VDDAI VSS TSMC_447 
+ TSMC_448 TSMC_319 TSMC_320 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD33 TSMC_61 TSMC_62 TSMC_189 TSMC_190 VSS VDDM VDDAI VSS TSMC_445 
+ TSMC_446 TSMC_317 TSMC_318 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD34 TSMC_59 TSMC_60 TSMC_187 TSMC_188 VSS VDDM VDDAI VSS TSMC_443 
+ TSMC_444 TSMC_315 TSMC_316 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD35 TSMC_57 TSMC_58 TSMC_185 TSMC_186 VSS VDDM VDDAI VSS TSMC_441 
+ TSMC_442 TSMC_313 TSMC_314 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD36 TSMC_55 TSMC_56 TSMC_183 TSMC_184 VSS VDDM VDDAI VSS TSMC_439 
+ TSMC_440 TSMC_311 TSMC_312 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD37 TSMC_53 TSMC_54 TSMC_181 TSMC_182 VSS VDDM VDDAI VSS TSMC_437 
+ TSMC_438 TSMC_309 TSMC_310 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD38 TSMC_51 TSMC_52 TSMC_179 TSMC_180 VSS VDDM VDDAI VSS TSMC_435 
+ TSMC_436 TSMC_307 TSMC_308 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD39 TSMC_49 TSMC_50 TSMC_177 TSMC_178 VSS VDDM VDDAI VSS TSMC_433 
+ TSMC_434 TSMC_305 TSMC_306 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD40 TSMC_47 TSMC_48 TSMC_175 TSMC_176 VSS VDDM VDDAI VSS TSMC_431 
+ TSMC_432 TSMC_303 TSMC_304 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD41 TSMC_45 TSMC_46 TSMC_173 TSMC_174 VSS VDDM VDDAI VSS TSMC_429 
+ TSMC_430 TSMC_301 TSMC_302 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD42 TSMC_43 TSMC_44 TSMC_171 TSMC_172 VSS VDDM VDDAI VSS TSMC_427 
+ TSMC_428 TSMC_299 TSMC_300 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD43 TSMC_41 TSMC_42 TSMC_169 TSMC_170 VSS VDDM VDDAI VSS TSMC_425 
+ TSMC_426 TSMC_297 TSMC_298 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD44 TSMC_39 TSMC_40 TSMC_167 TSMC_168 VSS VDDM VDDAI VSS TSMC_423 
+ TSMC_424 TSMC_295 TSMC_296 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD45 TSMC_37 TSMC_38 TSMC_165 TSMC_166 VSS VDDM VDDAI VSS TSMC_421 
+ TSMC_422 TSMC_293 TSMC_294 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD46 TSMC_35 TSMC_36 TSMC_163 TSMC_164 VSS VDDM VDDAI VSS TSMC_419 
+ TSMC_420 TSMC_291 TSMC_292 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD47 TSMC_33 TSMC_34 TSMC_161 TSMC_162 VSS VDDM VDDAI VSS TSMC_417 
+ TSMC_418 TSMC_289 TSMC_290 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD48 TSMC_31 TSMC_32 TSMC_159 TSMC_160 VSS VDDM VDDAI VSS TSMC_415 
+ TSMC_416 TSMC_287 TSMC_288 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD49 TSMC_29 TSMC_30 TSMC_157 TSMC_158 VSS VDDM VDDAI VSS TSMC_413 
+ TSMC_414 TSMC_285 TSMC_286 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD50 TSMC_27 TSMC_28 TSMC_155 TSMC_156 VSS VDDM VDDAI VSS TSMC_411 
+ TSMC_412 TSMC_283 TSMC_284 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD51 TSMC_25 TSMC_26 TSMC_153 TSMC_154 VSS VDDM VDDAI VSS TSMC_409 
+ TSMC_410 TSMC_281 TSMC_282 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD52 TSMC_23 TSMC_24 TSMC_151 TSMC_152 VSS VDDM VDDAI VSS TSMC_407 
+ TSMC_408 TSMC_279 TSMC_280 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD53 TSMC_21 TSMC_22 TSMC_149 TSMC_150 VSS VDDM VDDAI VSS TSMC_405 
+ TSMC_406 TSMC_277 TSMC_278 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD54 TSMC_19 TSMC_20 TSMC_147 TSMC_148 VSS VDDM VDDAI VSS TSMC_403 
+ TSMC_404 TSMC_275 TSMC_276 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD55 TSMC_17 TSMC_18 TSMC_145 TSMC_146 VSS VDDM VDDAI VSS TSMC_401 
+ TSMC_402 TSMC_273 TSMC_274 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD56 TSMC_15 TSMC_16 TSMC_143 TSMC_144 VSS VDDM VDDAI VSS TSMC_399 
+ TSMC_400 TSMC_271 TSMC_272 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD57 TSMC_13 TSMC_14 TSMC_141 TSMC_142 VSS VDDM VDDAI VSS TSMC_397 
+ TSMC_398 TSMC_269 TSMC_270 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD58 TSMC_11 TSMC_12 TSMC_139 TSMC_140 VSS VDDM VDDAI VSS TSMC_395 
+ TSMC_396 TSMC_267 TSMC_268 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD59 TSMC_9 TSMC_10 TSMC_137 TSMC_138 VSS VDDM VDDAI VSS TSMC_393 
+ TSMC_394 TSMC_265 TSMC_266 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD60 TSMC_7 TSMC_8 TSMC_135 TSMC_136 VSS VDDM VDDAI VSS TSMC_391 
+ TSMC_392 TSMC_263 TSMC_264 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD61 TSMC_5 TSMC_6 TSMC_133 TSMC_134 VSS VDDM VDDAI VSS TSMC_389 
+ TSMC_390 TSMC_261 TSMC_262 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD62 TSMC_3 TSMC_4 TSMC_131 TSMC_132 VSS VDDM VDDAI VSS TSMC_387 
+ TSMC_388 TSMC_259 TSMC_260 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLD63 TSMC_1 TSMC_2 TSMC_129 TSMC_130 VSS VDDM VDDAI VSS TSMC_385 
+ TSMC_386 TSMC_257 TSMC_258 TSMC_532 TSMC_533 TSMC_531 
+ S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X2 
XRWLLDL TSMC_513 TSMC_514 VSS VDDM VDDAI VSS TSMC_534 TSMC_515 TSMC_535 
+ TSMC_531 S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X1 
XRWLLDR TSMC_517 TSMC_514 VSS VDDM VDDAI VSS TSMC_536 TSMC_518 TSMC_535 
+ TSMC_531 S6ALLSVTFW40W20_D130_ARRAY_RWL_TRK_X1 
XDECCAP TSMC_537 TSMC_523 TSMC_520 TSMC_521 TSMC_522 VDDM VDDI VSS TSMC_515 
+ TSMC_519 TSMC_516 TSMC_524 TSMC_531 TSMC_531 
+ S6ALLSVTFW40W20_RF_XDECCAP 
.ENDS

.SUBCKT TS6N16FFCLLSVTA64X32M4FW D[31] D[30] D[29] D[28] D[27] D[26] D[25] 
+ D[24] D[23] D[22] D[21] D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] 
+ D[11] D[10] D[9] D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] Q[31] Q[30] 
+ Q[29] Q[28] Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] 
+ Q[16] Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] 
+ Q[2] Q[1] Q[0] BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] BWEB[25] 
+ BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] BWEB[18] BWEB[17] 
+ BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] BWEB[11] BWEB[10] BWEB[9] 
+ BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] BWEB[3] BWEB[2] BWEB[1] BWEB[0] AB[5] 
+ AB[4] AB[3] AB[2] AB[1] AB[0] CLKR REB AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] 
+ CLKW WEB KP[2] KP[1] KP[0] WCT[1] WCT[0] RCT[1] RCT[0] VDD VSS 
XPIN_ROW D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] D[22] D[21] 
+ D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] D[10] D[9] 
+ D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] Q[31] Q[30] Q[29] Q[28] 
+ Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] Q[16] 
+ Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] 
+ Q[2] Q[1] Q[0] BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] 
+ BWEB[25] BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] 
+ BWEB[18] BWEB[17] BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] 
+ BWEB[11] BWEB[10] BWEB[9] BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] 
+ BWEB[3] BWEB[2] BWEB[1] BWEB[0] TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] CLKR REB TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] CLKW WEB KP[2] KP[1] KP[0] 
+ TSMC_1 TSMC_2 TSMC_1 RCT[1] RCT[0] WCT[1] WCT[0] TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 VSS TSMC_3 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_2 TSMC_2 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_4 TSMC_5 TSMC_6 S6ALLSVTFW40W20_PIN_ROW 
XGCTRL_GIO CLKR CLKW D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] 
+ D[22] D[21] D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] 
+ D[10] D[9] D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 
+ TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 
+ TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 
+ TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 
+ TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 
+ TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 
+ TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 TSMC_155 
+ TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 
+ TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 KP[2] KP[1] KP[0] TSMC_168 
+ TSMC_169 TSMC_170 TSMC_1 TSMC_2 TSMC_1 TSMC_171 TSMC_172 TSMC_173 
+ TSMC_174 TSMC_175 TSMC_1 Q[31] Q[30] Q[29] Q[28] Q[27] Q[26] Q[25] 
+ Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] Q[16] Q[15] Q[14] Q[13] 
+ Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] 
+ RCT[1] RCT[0] REB TSMC_176 TSMC_1 TSMC_177 TSMC_178 TSMC_179 TSMC_180 
+ TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 
+ TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 
+ TSMC_195 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 AB[5] AB[4] AB[3] 
+ AB[2] TSMC_1 AB[1] AB[0] TSMC_1 TSMC_2 TSMC_1 TSMC_196 VDD VDD VSS 
+ TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 
+ TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 
+ TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 
+ TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 
+ TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 
+ TSMC_311 TSMC_312 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 
+ TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 
+ TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 
+ TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 
+ TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 
+ TSMC_375 TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 
+ TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 
+ TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 
+ TSMC_447 TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 WCT[1] WCT[0] WEB 
+ BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] BWEB[25] 
+ BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] BWEB[18] 
+ BWEB[17] BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] BWEB[11] 
+ BWEB[10] BWEB[9] BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] BWEB[3] 
+ BWEB[2] BWEB[1] BWEB[0] TSMC_453 TSMC_1 TSMC_454 TSMC_455 TSMC_456 
+ TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 
+ TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 
+ TSMC_472 TSMC_1 TSMC_1 TSMC_1 TSMC_1 AA[5] AA[4] AA[3] AA[2] TSMC_1 
+ AA[1] AA[0] TSMC_473 TSMC_1 TSMC_3 TSMC_474 TSMC_2 TSMC_475 TSMC_2 
+ TSMC_2 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 
+ TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 
+ TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 TSMC_525 
+ TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 TSMC_532 
+ TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 TSMC_539 TSMC_1 
+ S6ALLSVTFW40W20_GCTRL_GIO 
XROW_TRACKING TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 
+ TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 
+ TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 
+ TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 
+ TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 
+ TSMC_360 TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 
+ TSMC_367 TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 
+ TSMC_374 TSMC_375 TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 
+ TSMC_382 TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 
+ TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 
+ TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 
+ TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 
+ TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 
+ TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 
+ TSMC_425 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 
+ TSMC_432 TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 
+ TSMC_439 TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 
+ TSMC_447 TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_197 
+ TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 
+ TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 
+ TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 
+ TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 
+ TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 
+ TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 
+ TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 
+ TSMC_311 TSMC_312 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 
+ TSMC_318 TSMC_319 TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 
+ TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 
+ TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 
+ TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 
+ TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 
+ TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 
+ TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 
+ TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 VDD VDD VDD 
+ VSS TSMC_176 TSMC_176 TSMC_1 TSMC_196 TSMC_540 TSMC_541 
+ S6ALLSVTFW40W20_ROW_TRACKING 
XARY4ROW_SEG0_ARY0 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
+ TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 
+ TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 
+ TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 
+ TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 
+ TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 
+ TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 
+ TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 
+ TSMC_606 TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 
+ TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 
+ TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 
+ TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 
+ TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 
+ TSMC_664 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_325 
+ TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 
+ TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 
+ TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 
+ TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 
+ TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 
+ TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 
+ TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 
+ TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_670 TSMC_671 
+ TSMC_174 TSMC_167 TSMC_672 TSMC_673 TSMC_180 TSMC_181 TSMC_182 
+ TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 
+ TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_1 TSMC_1 VDD VDD 
+ VDD VSS TSMC_453 TSMC_454 TSMC_674 TSMC_457 TSMC_458 TSMC_459 TSMC_460 
+ TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_187 TSMC_191 
+ TSMC_464 TSMC_468 TSMC_540 TSMC_675 TSMC_541 TSMC_676 
+ TSMC_677 TSMC_678 TSMC_679 TSMC_680 S6ALLSVTFW40W20_ARY4ROW 
XARY4ROW_SEG0_ARY1 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
+ TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 
+ TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 
+ TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 
+ TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 
+ TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 
+ TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 
+ TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 
+ TSMC_606 TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 
+ TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 
+ TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 
+ TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 
+ TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 
+ TSMC_664 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_325 
+ TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 
+ TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 
+ TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 
+ TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 
+ TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 
+ TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 
+ TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 
+ TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_670 TSMC_671 
+ TSMC_174 TSMC_167 TSMC_672 TSMC_673 TSMC_180 TSMC_181 TSMC_182 
+ TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 
+ TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_1 TSMC_1 VDD VDD 
+ VDD VSS TSMC_453 TSMC_454 TSMC_674 TSMC_457 TSMC_458 TSMC_459 TSMC_460 
+ TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_186 TSMC_191 
+ TSMC_463 TSMC_468 TSMC_675 TSMC_681 TSMC_676 TSMC_682 
+ TSMC_678 TSMC_683 TSMC_680 TSMC_684 S6ALLSVTFW40W20_ARY4ROW 
XARY4ROW_SEG0_ARY2 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
+ TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 
+ TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 
+ TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 
+ TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 
+ TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 
+ TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 
+ TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 
+ TSMC_606 TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 
+ TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 
+ TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 
+ TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 
+ TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 
+ TSMC_664 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_325 
+ TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 
+ TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 
+ TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 
+ TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 
+ TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 
+ TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 
+ TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 
+ TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_670 TSMC_671 
+ TSMC_174 TSMC_167 TSMC_672 TSMC_673 TSMC_180 TSMC_181 TSMC_182 
+ TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 
+ TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_1 TSMC_1 VDD VDD 
+ VDD VSS TSMC_453 TSMC_454 TSMC_674 TSMC_457 TSMC_458 TSMC_459 TSMC_460 
+ TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_185 TSMC_191 
+ TSMC_462 TSMC_468 TSMC_681 TSMC_685 TSMC_682 TSMC_686 
+ TSMC_683 TSMC_687 TSMC_684 TSMC_688 S6ALLSVTFW40W20_ARY4ROW 
XARY4ROW_TK_SEG0_ARY3 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
+ TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 
+ TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 
+ TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 
+ TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 
+ TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 
+ TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 
+ TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 
+ TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 
+ TSMC_606 TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 
+ TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 
+ TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 
+ TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 
+ TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 
+ TSMC_664 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_325 
+ TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 
+ TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 
+ TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 
+ TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 
+ TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 
+ TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 
+ TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 
+ TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 
+ TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_670 TSMC_671 
+ TSMC_174 TSMC_167 TSMC_672 TSMC_673 TSMC_180 TSMC_181 TSMC_182 
+ TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 
+ TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_1 TSMC_1 VDD VDD 
+ VDD VSS TSMC_453 TSMC_454 TSMC_674 TSMC_457 TSMC_458 TSMC_459 TSMC_460 
+ TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_184 TSMC_191 
+ TSMC_461 TSMC_468 TSMC_685 TSMC_689 TSMC_686 TSMC_690 
+ TSMC_196 TSMC_196 TSMC_687 TSMC_691 TSMC_688 TSMC_692 
+ S6ALLSVTFW40W20_ARY4ROW_TK 
XLIO_LCTRL_SEG0 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 
+ TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_542 
+ TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 TSMC_561 
+ TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 TSMC_567 
+ TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 
+ TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 
+ TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 
+ TSMC_600 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 
+ TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 TSMC_612 
+ TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 
+ TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 TSMC_625 
+ TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 TSMC_631 
+ TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 
+ TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 TSMC_644 
+ TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 TSMC_657 
+ TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 TSMC_664 
+ TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_693 
+ TSMC_694 TSMC_695 TSMC_696 TSMC_697 TSMC_698 TSMC_699 TSMC_700 
+ TSMC_701 TSMC_702 TSMC_703 TSMC_704 TSMC_705 TSMC_706 
+ TSMC_707 TSMC_708 TSMC_709 TSMC_710 TSMC_711 TSMC_712 
+ TSMC_713 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 TSMC_719 
+ TSMC_720 TSMC_721 TSMC_722 TSMC_723 TSMC_724 TSMC_725 
+ TSMC_726 TSMC_727 TSMC_728 TSMC_729 TSMC_730 TSMC_731 TSMC_732 
+ TSMC_733 TSMC_734 TSMC_735 TSMC_736 TSMC_737 TSMC_738 
+ TSMC_739 TSMC_740 TSMC_741 TSMC_742 TSMC_743 TSMC_744 
+ TSMC_745 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 TSMC_751 
+ TSMC_752 TSMC_753 TSMC_754 TSMC_755 TSMC_756 TSMC_757 
+ TSMC_758 TSMC_759 TSMC_760 TSMC_761 TSMC_762 TSMC_763 TSMC_764 
+ TSMC_765 TSMC_766 TSMC_767 TSMC_768 TSMC_769 TSMC_770 
+ TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_775 TSMC_776 
+ TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_782 TSMC_783 
+ TSMC_784 TSMC_785 TSMC_786 TSMC_787 TSMC_788 TSMC_789 
+ TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_794 TSMC_795 TSMC_796 
+ TSMC_797 TSMC_798 TSMC_799 TSMC_800 TSMC_801 TSMC_802 
+ TSMC_803 TSMC_804 TSMC_805 TSMC_806 TSMC_807 TSMC_808 
+ TSMC_809 TSMC_810 TSMC_811 TSMC_812 TSMC_813 TSMC_814 TSMC_815 
+ TSMC_816 TSMC_817 TSMC_818 TSMC_819 TSMC_820 TSMC_325 TSMC_326 
+ TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 
+ TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 TSMC_340 
+ TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 TSMC_347 
+ TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 TSMC_355 
+ TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 TSMC_362 
+ TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 
+ TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 
+ TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 
+ TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 
+ TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 
+ TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 
+ TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 TSMC_412 
+ TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 TSMC_419 
+ TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 TSMC_426 TSMC_427 
+ TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 TSMC_434 
+ TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 TSMC_441 
+ TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 
+ TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_197 TSMC_198 TSMC_199 
+ TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 
+ TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 
+ TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 
+ TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 
+ TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 
+ TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 
+ TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 
+ TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 TSMC_298 TSMC_299 
+ TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 TSMC_306 
+ TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_821 TSMC_670 TSMC_821 
+ TSMC_1 TSMC_671 TSMC_176 TSMC_196 TSMC_1 TSMC_1 TSMC_1 TSMC_174 TSMC_175 
+ TSMC_196 TSMC_822 TSMC_167 TSMC_822 TSMC_196 TSMC_1 TSMC_1 TSMC_1 
+ VDD TSMC_473 TSMC_196 TSMC_191 TSMC_191 TSMC_168 TSMC_169 TSMC_170 
+ TSMC_171 TSMC_172 TSMC_173 TSMC_1 TSMC_823 TSMC_177 TSMC_673 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 
+ TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 
+ TSMC_195 TSMC_1 TSMC_1 TSMC_190 TSMC_190 VDD VDD VDD VSS TSMC_453 
+ TSMC_454 TSMC_674 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_176 TSMC_453 TSMC_824 TSMC_475 
+ TSMC_1 TSMC_825 TSMC_176 S6ALLSVTFW40W20_LIO_LCTRL 
XWRITE_TRAKING TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 
+ TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_542 
+ TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 TSMC_561 
+ TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 TSMC_567 
+ TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 
+ TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 
+ TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 
+ TSMC_600 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 
+ TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 TSMC_612 
+ TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 
+ TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 TSMC_625 
+ TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 TSMC_631 
+ TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 
+ TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 TSMC_644 
+ TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 TSMC_657 
+ TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 TSMC_664 
+ TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_197 
+ TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 
+ TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 
+ TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 
+ TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 
+ TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 
+ TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 
+ TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
+ TSMC_312 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 
+ TSMC_319 TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 
+ TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 
+ TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 
+ TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 
+ TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 
+ TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 
+ TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 TSMC_426 
+ TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 
+ TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_670 TSMC_671 TSMC_174 
+ TSMC_175 TSMC_167 TSMC_672 TSMC_473 TSMC_176 TSMC_823 TSMC_1 TSMC_1 
+ VDD VDD VDD VSS TSMC_453 TSMC_689 TSMC_690 TSMC_691 
+ TSMC_692 S6ALLSVTFW40W20_WRITE_TRAKING 
.ENDS


