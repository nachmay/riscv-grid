**** Created by MC2: Version 2013.12.00.f on 2025/06/22, 17:57:14 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  N16FF_SPSB_LEAFCELL
* Top Cell Name: LEAFCELL
* View Name:     schematic
* Netlisted on:  Jun  4 15:47:25 2014
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM


*.PIN vss
.SUBCKT ndio_mac PLUS MINUS 
.ends

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    XDRV_STRAP_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_XDRV_STRAP_SB TSMC_1 TSMC_2 VDDI VSSI 
MM10 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=6 m=20 
MM1 TSMC_2 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=3 m=10 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    BCELL_SD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_BCELL_SD TSMC_1 TSMC_2 VDDAI VDDI VSSI TSMC_3 
MM5 TSMC_2 TSMC_3 TSMC_4 VSSI nchpg_hcsr_mac l=20n nfin=2 m=1 
MM0 TSMC_1 TSMC_3 TSMC_5 VSSI nchpg_hcsr_mac l=20n nfin=2 m=1 
MM2 TSMC_4 TSMC_5 VSSI VSSI nchpd_hcsr_mac l=20n nfin=2 m=1 
MM1 TSMC_5 TSMC_4 VSSI VSSI nchpd_hcsr_mac l=20n nfin=2 m=1 
MM6 TSMC_5 TSMC_4 VDDAI VDDI pchpu_hcsr_mac l=20n nfin=1 m=1 
MM4 TSMC_4 TSMC_5 VDDAI VDDI pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_lvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_nand3_lvt_mac_pcell_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_lvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_lvt_mac_pcell_5
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_nor2_lvt_mac_pcell_5 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_6
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    XDRV_LA512_884_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_XDRV_LA512_884_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 VDDI VSSI TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 
MM37 TSMC_26 TSMC_30 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM36 TSMC_30 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM35 TSMC_22 TSMC_30 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM34 TSMC_30 TSMC_31 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM33 TSMC_31 TSMC_3 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MM21 TSMC_27 TSMC_33 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM16 TSMC_33 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM13 TSMC_23 TSMC_33 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM11 TSMC_33 TSMC_34 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM10 TSMC_34 TSMC_4 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MM3 TSMC_25 TSMC_35 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM2 TSMC_24 TSMC_36 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM23 TSMC_21 TSMC_35 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM20 TSMC_20 TSMC_36 VDDI VDDI pch_svt_mac l=20n nfin=8 m=8 
MM28 TSMC_35 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM27 TSMC_36 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM26 TSMC_35 TSMC_37 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM18 TSMC_36 TSMC_38 VDDI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM12 TSMC_37 TSMC_2 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MP6 TSMC_38 TSMC_1 TSMC_32 VDDI pch_svt_mac l=20n nfin=7 m=1 
MM39 TSMC_32 TSMC_9 VDDI VDDI pch_svt_mac l=20n nfin=7 m=4 
MM32 TSMC_26 TSMC_30 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM31 TSMC_22 TSMC_30 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM30 TSMC_30 TSMC_31 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM29 TSMC_31 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM22 TSMC_31 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM9 TSMC_27 TSMC_33 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM8 TSMC_23 TSMC_33 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM7 TSMC_33 TSMC_34 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM5 TSMC_34 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_34 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_25 TSMC_35 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM0 TSMC_24 TSMC_36 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM24 TSMC_21 TSMC_35 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM19 TSMC_20 TSMC_36 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM25 TSMC_35 TSMC_37 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM17 TSMC_36 TSMC_38 TSMC_29 VSSI nch_svt_mac l=20n nfin=12 m=1 
MM14 TSMC_37 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM6 TSMC_38 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM15 TSMC_37 TSMC_2 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MP9 TSMC_38 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    PRECHARGE_SB_SD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_PRECHARGE_SB_SD TSMC_1 TSMC_2 TSMC_3 VDDAI VDDI 
MM0_HDM VDDAI TSMC_3 TSMC_1 VDDI pch_svt_mac l=20n nfin=5 m=2 
MP5_HDM TSMC_1 TSMC_3 TSMC_2 VDDI pch_svt_mac l=20n nfin=5 m=1 
MP17_HDM TSMC_2 TSMC_3 VDDAI VDDI pch_svt_mac l=20n nfin=5 m=2 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MCB_2X4_SD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_MCB_2X4_SD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDAI VDDI VSSI TSMC_9 TSMC_10 
XMCB_0<0> TSMC_1 TSMC_5 VDDAI VDDI VSSI TSMC_9 
+ S1ALLSVTSW400W20_BCELL_SD 
XMCB_0<1> TSMC_2 TSMC_6 VDDAI VDDI VSSI TSMC_9 
+ S1ALLSVTSW400W20_BCELL_SD 
XMCB_0<2> TSMC_3 TSMC_7 VDDAI VDDI VSSI TSMC_9 
+ S1ALLSVTSW400W20_BCELL_SD 
XMCB_0<3> TSMC_4 TSMC_8 VDDAI VDDI VSSI TSMC_9 
+ S1ALLSVTSW400W20_BCELL_SD 
XMCB_1<0> TSMC_1 TSMC_5 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW400W20_BCELL_SD 
XMCB_1<1> TSMC_2 TSMC_6 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW400W20_BCELL_SD 
XMCB_1<2> TSMC_3 TSMC_7 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW400W20_BCELL_SD 
XMCB_1<3> TSMC_4 TSMC_8 VDDAI VDDI VSSI TSMC_10 
+ S1ALLSVTSW400W20_BCELL_SD 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MIO_M4_SB_BUF
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_MIO_M4_SB_BUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VSSI 
XI8 VSSI VSSI TSMC_6 TSMC_7 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI9 VSSI VSSI TSMC_7 TSMC_4 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI15 VSSI VSSI TSMC_8 TSMC_2 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI14 VSSI VSSI TSMC_9 TSMC_8 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI16 VSSI VSSI TSMC_3 TSMC_6 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI17 VSSI VSSI TSMC_1 TSMC_9 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DIO_TALL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DIO_TALL TSMC_1 TSMC_2 
XDDIO_TALL TSMC_2 TSMC_1 ndio_mac nfin=2 l=2e-07 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    XDRV_STRAP_BT_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_XDRV_STRAP_BT_SB TSMC_1 TSMC_2 VDDI VSSI 
MM0 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=12 m=4 
MM10 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=6 m=12 
MM1 TSMC_2 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=3 m=10 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    RESETD_WTSEL_SB_NEW
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_RESETD_WTSEL_SB_NEW TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ TSMC_3 TSMC_4 
XI87 TSMC_5 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_7 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND5 TSMC_4 TSMC_8 VSSI VSSI VDDHD VDDI TSMC_5 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI84 TSMC_3 TSMC_9 VSSI VSSI VDDHD VDDI TSMC_6 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND0 TSMC_5 TSMC_1 VSSI VSSI VDDHD VDDI TSMC_9 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI89 VSSI VSSI TSMC_7 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI65 VSSI VSSI TSMC_10 TSMC_11 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI83 VSSI VSSI TSMC_11 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI64 VSSI VSSI TSMC_1 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    RESETD_TSEL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_RESETD_TSEL TSMC_1 TSMC_2 TSMC_3 VDDHD VDDI VSSI 
+ TSMC_4 TSMC_5 
MM15 TSMC_6 TSMC_1 TSMC_7 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14 TSMC_7 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM25 TSMC_4 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM23 TSMC_4 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM18 TSMC_6 TSMC_1 TSMC_9 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM19 TSMC_9 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM24 TSMC_10 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM21 TSMC_4 TSMC_2 TSMC_10 VSSI nch_svt_mac l=20n nfin=3 m=1 
XI737 VSSI VSSI TSMC_11 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI736 VSSI VSSI TSMC_12 TSMC_11 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XND0 TSMC_1 TSMC_5 VSSI VSSI VDDHD VDDI TSMC_8 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI91 TSMC_3 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_12 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    WEBBUF_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_WEBBUF_SB_BASE TSMC_1 TSMC_2 VDDHD VDDI VSSI TSMC_3 
+ TSMC_4 TSMC_5 
MM36 TSMC_6 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM35 TSMC_8 TSMC_2 TSMC_6 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM31 TSMC_9 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=5 m=2 
MM30 TSMC_8 TSMC_3 TSMC_9 VSSI nch_svt_mac l=20n nfin=5 m=1 
MM34 TSMC_10 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM33 TSMC_8 TSMC_1 TSMC_10 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM6 TSMC_8 TSMC_3 TSMC_11 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM32 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
XI25 VSSI VSSI TSMC_8 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI32 VSSI VSSI TSMC_8 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=7 p_l=20n 
XI33 VSSI VSSI TSMC_5 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB4_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 VDDHD VDDI VSSI 
MM15 TSMC_10 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM16 TSMC_10 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM17 TSMC_11 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM18 TSMC_11 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM22 TSMC_11 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM23 TSMC_10 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM24 TSMC_12 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM25 TSMC_13 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_12 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_12 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM2 TSMC_13 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_13 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM19 TSMC_14 TSMC_4 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=2 
MM20 TSMC_10 TSMC_2 TSMC_14 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM21 TSMC_11 TSMC_1 TSMC_14 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM26 TSMC_15 TSMC_5 VSSI VSSI nch_svt_mac l=20n nfin=3 m=4 
MM8 TSMC_16 TSMC_3 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=2 
MM7 TSMC_12 TSMC_2 TSMC_16 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM0 TSMC_13 TSMC_1 TSMC_16 VSSI nch_svt_mac l=20n nfin=3 m=1 
XINV3 VSSI VSSI TSMC_10 TSMC_9 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV2 VSSI VSSI TSMC_11 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV1 VSSI VSSI TSMC_12 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV0 VSSI VSSI TSMC_13 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB1_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VDDHD VDDI VSSI 
MTN1 TSMC_8 TSMC_1 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_9 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MM0 TSMC_8 TSMC_2 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=4 
MM1 TSMC_10 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_8 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=6 
MP5 TSMC_8 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_8 TSMC_1 TSMC_10 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB2_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB2_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD VDDI 
+ VSSI 
MM2 TSMC_6 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_6 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_7 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_7 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM0 TSMC_6 TSMC_1 TSMC_8 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_7 TSMC_2 TSMC_8 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM8 TSMC_8 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=3 m=2 
XINV0 VSSI VSSI TSMC_7 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XINV1 VSSI VSSI TSMC_6 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_BLEQ_SB_M4
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB1_BLEQ_SB_M4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 VDDHD VDDI VSSI 
MN0 TSMC_1 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=8 m=4 
MTN1 TSMC_7 TSMC_3 TSMC_6 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MM0 TSMC_7 TSMC_4 TSMC_6 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM2 TSMC_2 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=8 m=4 
MP0 TSMC_1 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=6 
MM4 TSMC_7 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM3 TSMC_7 TSMC_3 TSMC_8 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_8 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_2 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=6 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_WLNAD2_SB_X0
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD VDDI VSSI 
MM5 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MTN1 TSMC_9 TSMC_1 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_10 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM0 TSMC_9 TSMC_2 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=6 
MM4 TSMC_8 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MM1 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_9 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=3 
MP5 TSMC_9 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CKBUF_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_CKBUF_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI VSSI 
XINV0 VSSI VSSI TSMC_1 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=7 n_l=20n p_totalM=3 
+ p_nfin=9 p_l=20n 
MM1 TSMC_1 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM34 TSMC_1 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=7 m=2 
MM26 TSMC_5 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=9 m=2 
MM0 TSMC_1 TSMC_4 TSMC_5 VDDI pch_svt_mac l=20n nfin=9 m=2 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    ABUF_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_ABUF_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VSSI 
MM15 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM14 TSMC_3 TSMC_5 TSMC_8 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM9 TSMC_10 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM8 TSMC_3 TSMC_1 TSMC_10 VSSI nch_svt_mac l=20n nfin=4 m=1 
MM13 TSMC_11 TSMC_9 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM12 TSMC_3 TSMC_4 TSMC_11 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM11 TSMC_3 TSMC_1 TSMC_12 TSMC_6 pch_svt_mac l=20n nfin=5 m=1 
MM10 TSMC_12 TSMC_5 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=5 m=2 
XI34 VSSI VSSI TSMC_3 TSMC_9 TSMC_7 TSMC_6 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI35 VSSI VSSI TSMC_3 TSMC_2 TSMC_7 TSMC_6 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    ENBUFB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_ENBUFB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDHD VDDI VSSI 
XI158 TSMC_9 TSMC_9 VSSI VSSI VDDHD VDDI TSMC_10 
+ S1ALLSVTSW400W20_nor2_lvt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM19 TSMC_11 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=6 m=1 
MM2 TSMC_12 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_13 TSMC_8 VDDI VDDI pch_svt_mac l=20n nfin=5 m=1 
MM16 TSMC_13 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=6 m=1 
MM1 TSMC_13 TSMC_2 TSMC_12 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_14 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN200 TSMC_6 TSMC_4 VSSI VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MM4 TSMC_15 TSMC_4 TSMC_14 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_13 TSMC_3 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM20 TSMC_16 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=7 m=1 
MM17 TSMC_13 TSMC_1 TSMC_17 VSSI nch_svt_mac l=20n nfin=4 m=1 
MM18 TSMC_17 TSMC_2 TSMC_16 VSSI nch_svt_mac l=20n nfin=4 m=1 
MN300 TSMC_5 TSMC_4 VSSI VSSI nch_ulvt_mac l=20n nfin=11 m=6 
XI166 VSSI VSSI TSMC_18 TSMC_9 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI148 VSSI VSSI TSMC_4 TSMC_18 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI152 VSSI VSSI TSMC_19 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=4 n_nfin=4 n_l=20n p_totalM=4 
+ p_nfin=8 p_l=20n 
XINV5 VSSI VSSI TSMC_4 TSMC_19 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=3 
+ p_nfin=3 p_l=20n 
XINV4 VSSI VSSI TSMC_10 TSMC_20 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI141 VSSI VSSI TSMC_13 TSMC_4 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=7 n_l=20n p_totalM=3 
+ p_nfin=9 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_WLNAD2_SB_X1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD VDDI VSSI 
MM5 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MTN1 TSMC_9 TSMC_1 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_10 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM0 TSMC_9 TSMC_2 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=6 
MM4 TSMC_8 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MM1 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_9 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=3 
MP5 TSMC_9 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MIO_SB_EDGE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_MIO_SB_EDGE VDDI TSMC_1 TSMC_2 VSSI 
MP0 TSMC_3 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP2 TSMC_4 TSMC_5 VDDI VDDI pch_svt_mac l=20n nfin=3 m=6 
MP7 TSMC_3 TSMC_5 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MN3 VSSI TSMC_3 TSMC_5 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1 VSSI TSMC_3 TSMC_6 VSSI nch_svt_mac l=20n nfin=3 m=5 
MN0 VSSI TSMC_5 TSMC_5 VSSI nch_svt_mac l=20n nfin=3 m=1 
XI18 VSSI VSSI TSMC_4 TSMC_2 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=8 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI393 VSSI VSSI TSMC_6 TSMC_1 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=4 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CKG_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_CKG_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD VDDI 
+ VSSI 
XI58 VSSI VSSI TSMC_6 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM0 TSMC_1 TSMC_7 VDDHD VDDI pch_svt_mac l=16.0n nfin=4 m=1 
MM26 TSMC_1 TSMC_8 VDDHD VDDI pch_svt_mac l=16.0n nfin=4 m=4 
MM1 TSMC_9 TSMC_8 VSSI VSSI nch_svt_mac l=16.0n nfin=8 m=3 
MM34 TSMC_1 TSMC_7 TSMC_9 VSSI nch_svt_mac l=16.0n nfin=8 m=3 
XNAND2 TSMC_2 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_10 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND5 TSMC_4 TSMC_1 VSSI VSSI VDDI VDDI TSMC_7 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND0 TSMC_1 TSMC_5 VSSI VSSI VDDHD VDDI TSMC_11 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND3 TSMC_10 TSMC_11 VSSI VSSI VDDHD VDDI TSMC_6 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XNAND12 TSMC_2 TSMC_3 TSMC_4 VSSI VSSI VDDI VDDI TSMC_8 
+ S1ALLSVTSW400W20_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=10 n_l=16.0n 
+ p_totalM=1 p_nfin=4 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    RESETD_884_M4_SB_NBL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_RESETD_884_M4_SB_NBL TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDDHD VDDI VSSI TSMC_12 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
XTSEL_WT TSMC_19 TSMC_20 VDDHD VDDI VSSI TSMC_16 TSMC_17 
+ S1ALLSVTSW400W20_RESETD_WTSEL_SB_NEW 
MM10 TSMC_21 TSMC_9 TSMC_11 VDDI pch_svt_mac l=16.0n nfin=3 m=1 
MP0 TSMC_11 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=4 m=3 
MM0 TSMC_22 TSMC_23 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MI537 TSMC_1 TSMC_23 VDDHD VDDI pch_svt_mac l=16.0n nfin=8 m=4 
MM5 TSMC_21 TSMC_24 TSMC_25 VDDI pch_svt_mac l=20n nfin=3 m=1 
XTSEL_READ TSMC_3 TSMC_14 TSMC_15 VDDHD VDDI VSSI TSMC_26 TSMC_27 
+ S1ALLSVTSW400W20_RESETD_TSEL 
MM12 TSMC_21 TSMC_24 TSMC_11 VSSI nch_svt_mac l=16.0n nfin=4 m=2 
MM11 TSMC_1 TSMC_23 VSSI VSSI nch_svt_mac l=16.0n nfin=5 m=4 
MM4 TSMC_21 TSMC_9 TSMC_25 VSSI nch_svt_mac l=20n nfin=4 m=2 
MM1 TSMC_8 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=5 m=1 
XNAND3 TSMC_27 TSMC_26 TSMC_3 VSSI VSSI VDDI VDDI TSMC_23 
+ S1ALLSVTSW400W20_nand3_lvt_mac_pcell_2 n_totalM=2 n_nfin=9 n_l=16.0n 
+ p_totalM=2 p_nfin=3 p_l=16.0n 
XI667 TSMC_19 TSMC_2 TSMC_28 VSSI VSSI VDDHD VDDI TSMC_29 
+ S1ALLSVTSW400W20_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=9 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XI696 TSMC_19 TSMC_20 VSSI VSSI VDDHD VDDI TSMC_30 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI658 TSMC_18 TSMC_1 VSSI VSSI VDDHD VDDI TSMC_31 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI728 TSMC_1 TSMC_32 VSSI VSSI VDDHD VDDI TSMC_25 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI666 TSMC_29 TSMC_33 VSSI VSSI VDDHD VDDI TSMC_34 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XI654 TSMC_31 TSMC_30 VSSI VSSI TSMC_22 VDDI TSMC_8 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI725 VSSI VSSI TSMC_9 TSMC_24 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI730 VSSI VSSI TSMC_35 TSMC_36 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI731 VSSI VSSI TSMC_36 TSMC_37 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI732 VSSI VSSI TSMC_37 TSMC_38 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI733 VSSI VSSI TSMC_38 TSMC_28 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI703 VSSI VSSI TSMC_12 TSMC_35 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI695 VSSI VSSI TSMC_39 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=3 n_nfin=6 n_l=20n p_totalM=4 
+ p_nfin=7 p_l=20n 
XI679 VSSI VSSI TSMC_34 TSMC_40 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=9 n_l=16.0n p_totalM=1 
+ p_nfin=8 p_l=16.0n 
XI693 VSSI VSSI TSMC_3 TSMC_39 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XI713 VSSI VSSI TSMC_21 TSMC_19 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=16.0n p_totalM=2 
+ p_nfin=3 p_l=16.0n 
XI718 VSSI VSSI TSMC_6 TSMC_32 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI686 VSSI VSSI TSMC_41 TSMC_33 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI687 VSSI VSSI TSMC_40 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=8 n_nfin=7 n_l=16.0n p_totalM=8 
+ p_nfin=10 p_l=16.0n 
XI685 VSSI VSSI TSMC_31 TSMC_41 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    COTH_M4_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_COTH_M4_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ VSSI TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
XCKG TSMC_5 TSMC_7 TSMC_8 TSMC_9 TSMC_25 TSMC_16 TSMC_15 VSSI 
+ S1ALLSVTSW400W20_CKG_SB 
XWEBBUF TSMC_3 TSMC_4 TSMC_16 TSMC_15 VSSI TSMC_17 TSMC_18 TSMC_19 
+ S1ALLSVTSW400W20_WEBBUF_SB_BASE 
XRESETD TSMC_1 TSMC_2 TSMC_5 TSMC_6 TSMC_26 TSMC_7 TSMC_21 TSMC_25 TSMC_12 
+ TSMC_13 TSMC_14 TSMC_16 TSMC_15 VSSI TSMC_19 TSMC_20 TSMC_10 TSMC_11 
+ TSMC_22 TSMC_23 TSMC_24 S1ALLSVTSW400W20_RESETD_884_M4_SB_NBL 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_Y_M4_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB1_Y_M4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD VDDI VSSI 
MM6 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=9 m=9 
MTN1 TSMC_9 TSMC_1 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_10 TSMC_7 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM0 TSMC_9 TSMC_2 TSMC_10 VSSI nch_ulvt_mac l=20n nfin=6 m=2 
MM7 TSMC_8 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=7 m=6 
MM3 TSMC_9 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP5 TSMC_9 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM1 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM2 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DECB1_DCLK_M4_SB_V2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DECB1_DCLK_M4_SB_V2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 VDDHD VDDI VSSI 
MM2 TSMC_4 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=5 
MTN1 TSMC_8 TSMC_1 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_9 TSMC_7 TSMC_6 VSSI nch_ulvt_mac l=20n nfin=6 m=4 
MM0 TSMC_8 TSMC_2 TSMC_9 VSSI nch_ulvt_mac l=20n nfin=6 m=4 
MN0 TSMC_3 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=8 m=5 
MM4 TSMC_4 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=8 
MM1 TSMC_10 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_8 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=8 m=8 
MP5 TSMC_8 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=2 
MM5 TSMC_8 TSMC_1 TSMC_10 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CDEC_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_CDEC_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 VSSI TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 
XPREDEC_Y<0> TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_47 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_45 TSMC_44 VSSI S1ALLSVTSW400W20_DECB4_SB 
XPREDEC_Y<1> TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_48 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_45 TSMC_44 VSSI S1ALLSVTSW400W20_DECB4_SB 
XIPDEC_X1<0> TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 
+ TSMC_83 TSMC_45 TSMC_44 VSSI S1ALLSVTSW400W20_DECB4_SB 
XIPDEC_X1<1> TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_45 TSMC_44 VSSI S1ALLSVTSW400W20_DECB4_SB 
XIPDEC_X0<0> TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_45 TSMC_44 VSSI S1ALLSVTSW400W20_DECB4_SB 
XIPDEC_X0<1> TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_98 TSMC_99 TSMC_100 TSMC_101 
+ TSMC_102 TSMC_45 TSMC_44 VSSI S1ALLSVTSW400W20_DECB4_SB 
XIDEC_X2<0> TSMC_8 TSMC_10 TSMC_28 TSMC_40 TSMC_103 TSMC_41 TSMC_104 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_SB 
XIDEC_X2<1> TSMC_8 TSMC_10 TSMC_29 TSMC_40 TSMC_103 TSMC_41 TSMC_105 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_SB 
XIDEC_X2<2> TSMC_8 TSMC_10 TSMC_30 TSMC_40 TSMC_103 TSMC_41 TSMC_106 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_SB 
XIDEC_X2<3> TSMC_8 TSMC_10 TSMC_31 TSMC_40 TSMC_103 TSMC_41 TSMC_107 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_SB 
XI381<0> TSMC_108 TSMC_109 TSMC_110 TSMC_104 TSMC_105 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW400W20_DECB2_SB 
XI381<1> TSMC_108 TSMC_109 TSMC_111 TSMC_106 TSMC_107 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW400W20_DECB2_SB 
XDECB1_BLEQ TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_112 TSMC_113 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW400W20_DECB1_BLEQ_SB_M4 
XIDEC_X0<0> TSMC_9 TSMC_10 TSMC_12 TSMC_112 TSMC_113 TSMC_41 TSMC_94 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XIDEC_X0<1> TSMC_9 TSMC_10 TSMC_13 TSMC_112 TSMC_113 TSMC_41 TSMC_95 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XIDEC_X0<2> TSMC_9 TSMC_10 TSMC_14 TSMC_112 TSMC_113 TSMC_41 TSMC_96 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XIDEC_X0<3> TSMC_9 TSMC_10 TSMC_15 TSMC_112 TSMC_113 TSMC_41 TSMC_97 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XIDEC_X0<4> TSMC_9 TSMC_10 TSMC_16 TSMC_112 TSMC_113 TSMC_41 TSMC_99 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XIDEC_X0<5> TSMC_9 TSMC_10 TSMC_17 TSMC_112 TSMC_113 TSMC_41 TSMC_100 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XIDEC_X0<6> TSMC_9 TSMC_10 TSMC_18 TSMC_112 TSMC_113 TSMC_41 TSMC_101 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XIDEC_X0<7> TSMC_9 TSMC_10 TSMC_19 TSMC_112 TSMC_113 TSMC_41 TSMC_102 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X0 
XCKBUF TSMC_4 TSMC_5 TSMC_9 TSMC_11 TSMC_45 TSMC_44 VSSI 
+ S1ALLSVTSW400W20_CKBUF_SB 
XABUF_Y<0> TSMC_57 TSMC_63 TSMC_64 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_Y<1> TSMC_58 TSMC_65 TSMC_66 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<3> TSMC_52 TSMC_75 TSMC_76 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<4> TSMC_53 TSMC_77 TSMC_78 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<5> TSMC_54 TSMC_79 TSMC_84 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<6> TSMC_55 TSMC_108 TSMC_109 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<7> TSMC_56 TSMC_110 TSMC_111 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<0> TSMC_49 TSMC_89 TSMC_90 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<1> TSMC_50 TSMC_91 TSMC_92 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XABUF_X<2> TSMC_51 TSMC_93 TSMC_98 TSMC_4 TSMC_5 TSMC_44 TSMC_45 VSSI 
+ S1ALLSVTSW400W20_ABUF_SB_BASE 
XIDEC_Y<0> TSMC_9 TSMC_10 TSMC_32 TSMC_112 TSMC_113 TSMC_41 TSMC_67 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_Y<1> TSMC_9 TSMC_10 TSMC_33 TSMC_112 TSMC_113 TSMC_41 TSMC_68 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_Y<2> TSMC_9 TSMC_10 TSMC_34 TSMC_112 TSMC_113 TSMC_41 TSMC_69 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_Y<3> TSMC_9 TSMC_10 TSMC_35 TSMC_112 TSMC_113 TSMC_41 TSMC_70 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_Y<4> TSMC_9 TSMC_11 TSMC_36 TSMC_112 TSMC_113 TSMC_41 TSMC_71 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_Y<5> TSMC_9 TSMC_11 TSMC_37 TSMC_112 TSMC_113 TSMC_41 TSMC_72 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_Y<6> TSMC_9 TSMC_11 TSMC_38 TSMC_112 TSMC_113 TSMC_41 TSMC_73 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_Y<7> TSMC_9 TSMC_11 TSMC_39 TSMC_112 TSMC_113 TSMC_41 TSMC_74 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_Y_M4_SB 
XIDEC_CKD TSMC_9 TSMC_10 TSMC_6 TSMC_7 TSMC_112 TSMC_113 TSMC_48 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_DCLK_M4_SB_V2 
XIDEC_X1<0> TSMC_9 TSMC_10 TSMC_20 TSMC_112 TSMC_113 TSMC_41 TSMC_80 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XIDEC_X1<1> TSMC_9 TSMC_10 TSMC_21 TSMC_112 TSMC_113 TSMC_41 TSMC_81 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XIDEC_X1<2> TSMC_9 TSMC_10 TSMC_22 TSMC_112 TSMC_113 TSMC_41 TSMC_82 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XIDEC_X1<3> TSMC_9 TSMC_10 TSMC_23 TSMC_112 TSMC_113 TSMC_41 TSMC_83 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XIDEC_X1<4> TSMC_9 TSMC_10 TSMC_24 TSMC_112 TSMC_113 TSMC_41 TSMC_85 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XIDEC_X1<5> TSMC_9 TSMC_10 TSMC_25 TSMC_112 TSMC_113 TSMC_41 TSMC_86 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XIDEC_X1<6> TSMC_9 TSMC_10 TSMC_26 TSMC_112 TSMC_113 TSMC_41 TSMC_87 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XIDEC_X1<7> TSMC_9 TSMC_10 TSMC_27 TSMC_112 TSMC_113 TSMC_41 TSMC_88 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_DECB1_WLNAD2_SB_X1 
XCEBBUF TSMC_3 TSMC_4 TSMC_5 TSMC_40 TSMC_113 TSMC_103 TSMC_112 TSMC_43 TSMC_45 
+ TSMC_44 VSSI S1ALLSVTSW400W20_ENBUFB_BASE 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CNT_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_CNT_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 VSSI TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 
XCOTHERS TSMC_3 TSMC_3 TSMC_65 TSMC_66 TSMC_7 TSMC_67 TSMC_8 TSMC_68 TSMC_69 
+ TSMC_42 TSMC_43 TSMC_45 TSMC_70 TSMC_46 TSMC_47 TSMC_47 VSSI TSMC_48 
+ TSMC_71 TSMC_49 TSMC_44 TSMC_72 TSMC_50 TSMC_51 TSMC_52 
+ S1ALLSVTSW400W20_COTH_M4_BASE 
Xcdec TSMC_1 TSMC_2 TSMC_4 TSMC_65 TSMC_66 TSMC_5 TSMC_6 TSMC_7 TSMC_67 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_68 TSMC_73 TSMC_74 
+ TSMC_69 TSMC_47 TSMC_47 VSSI TSMC_75 TSMC_71 TSMC_49 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_76 TSMC_77 S1ALLSVTSW400W20_CDEC_M4_SB_BASE 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DIN_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DIN_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI 
+ VSSI TSMC_5 TSMC_6 
MM6 TSMC_7 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM4 TSMC_9 TSMC_10 TSMC_11 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM35 TSMC_12 TSMC_13 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM41 TSMC_14 TSMC_13 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN33 TSMC_7 TSMC_15 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM19 TSMC_16 TSMC_1 TSMC_17 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM1 VSSI TSMC_8 TSMC_18 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM12 TSMC_16 TSMC_10 TSMC_14 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM5 VSSI TSMC_19 TSMC_11 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM9 TSMC_20 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM42 TSMC_17 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM34 TSMC_9 TSMC_3 TSMC_18 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM8 TSMC_20 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=2 m=2 
MM39 TSMC_22 TSMC_10 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM26 VDDHD TSMC_10 TSMC_23 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_24 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=4 
MM2 VDDHD TSMC_19 TSMC_25 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM33 TSMC_21 TSMC_13 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM36 TSMC_15 TSMC_13 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_9 TSMC_8 TSMC_25 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM14 TSMC_20 TSMC_21 TSMC_24 VDDI pch_svt_mac l=20n nfin=3 m=2 
MM0 TSMC_9 TSMC_3 TSMC_23 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM51 TSMC_7 TSMC_15 TSMC_24 VDDI pch_svt_mac l=20n nfin=3 m=2 
MM16 TSMC_16 TSMC_8 TSMC_26 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM15 TSMC_16 TSMC_1 TSMC_22 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM40 TSMC_26 TSMC_13 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
XI395 TSMC_12 VSSI TSMC_9 TSMC_21 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI295 TSMC_4 VSSI TSMC_7 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=3 n_nfin=9 n_l=20n p_totalM=3 
+ p_nfin=2 p_l=20n 
XI341 VSSI VSSI TSMC_2 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI396 TSMC_12 VSSI TSMC_19 TSMC_15 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI277 VSSI VSSI TSMC_16 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI339 TSMC_4 VSSI TSMC_20 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=3 n_nfin=9 n_l=20n p_totalM=3 
+ p_nfin=2 p_l=20n 
XI386 VSSI VSSI TSMC_8 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XINV04 VSSI VSSI TSMC_9 TSMC_19 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DOUT_SB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DOUT_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD VDDI 
+ VSSI 
MP11 TSMC_6 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM12 TSMC_6 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM9 TSMC_8 TSMC_7 TSMC_6 VDDI pch_svt_mac l=20n nfin=5 m=2 
MM17 TSMC_9 TSMC_10 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM8 TSMC_8 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MP14 TSMC_6 TSMC_12 TSMC_3 VDDI pch_svt_mac l=20n nfin=5 m=1 
MP13 TSMC_8 TSMC_12 TSMC_2 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM14_SA TSMC_13 TSMC_8 VDDHD VDDI pch_lvt_mac l=20n nfin=6 m=1 
MP2 TSMC_8 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MP10 TSMC_4 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=4 m=4 
MM35_SA TSMC_14 TSMC_6 VDDHD VDDI pch_lvt_mac l=20n nfin=6 m=1 
MM24_SA TSMC_15 TSMC_16 TSMC_14 VDDI pch_lvt_mac l=20n nfin=6 m=1 
MM20 TSMC_11 TSMC_17 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM23_SA TSMC_9 TSMC_16 TSMC_13 VDDI pch_lvt_mac l=20n nfin=6 m=1 
MM31_SA TSMC_18 TSMC_6 VSSI VSSI nch_lvt_mac l=20n nfin=3 m=1 
MN1 TSMC_6 TSMC_8 TSMC_19 VSSI nch_svt_mac l=20n nfin=10 m=4 
MM7 TSMC_19 TSMC_10 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM6 TSMC_8 TSMC_6 TSMC_19 VSSI nch_svt_mac l=20n nfin=10 m=4 
MM15_SA TSMC_20 TSMC_8 VSSI VSSI nch_lvt_mac l=20n nfin=3 m=1 
MM13_SA TSMC_9 TSMC_10 TSMC_20 VSSI nch_lvt_mac l=20n nfin=3 m=1 
MM18 TSMC_9 TSMC_16 TSMC_21 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN5 TSMC_4 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=4 m=4 
MM29_SA TSMC_15 TSMC_10 TSMC_18 VSSI nch_lvt_mac l=20n nfin=3 m=1 
MM21 TSMC_21 TSMC_17 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
XIPGB0 TSMC_22 TSMC_16 TSMC_7 VSSI VSSI VDDHD VDDI TSMC_12 
+ S1ALLSVTSW400W20_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI159 TSMC_16 TSMC_23 VSSI VSSI VDDHD VDDI TSMC_7 
+ S1ALLSVTSW400W20_nand2_lvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI185 VSSI VSSI TSMC_16 TSMC_24 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI203 VSSI VSSI TSMC_25 TSMC_23 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI184 VSSI VSSI TSMC_10 TSMC_16 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI161 VSSI VSSI TSMC_26 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI194 VSSI VSSI TSMC_5 TSMC_26 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI186 VSSI VSSI TSMC_24 TSMC_22 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI201 VSSI VSSI TSMC_1 TSMC_25 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI163 VSSI VSSI TSMC_9 TSMC_17 VDDHD VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    YPASS_M4_SB_NBL_V2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_YPASS_M4_SB_NBL_V2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 VDDI VSSI TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
XI250<4> TSMC_13 VSSI TSMC_20 TSMC_24 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI250<5> TSMC_13 VSSI TSMC_21 TSMC_25 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI250<6> TSMC_13 VSSI TSMC_22 TSMC_26 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI250<7> TSMC_13 VSSI TSMC_23 TSMC_27 VDDI VDDI 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MN18<0> TSMC_5 TSMC_24 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN18<1> TSMC_6 TSMC_25 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN18<2> TSMC_7 TSMC_26 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN18<3> TSMC_8 TSMC_27 TSMC_14 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<0> TSMC_1 TSMC_24 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<1> TSMC_2 TSMC_25 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<2> TSMC_3 TSMC_26 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MN31<3> TSMC_4 TSMC_27 TSMC_15 VSSI nch_ulvt_mac l=20n nfin=7 m=2 
MM4 TSMC_10 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM0 TSMC_28 TSMC_10 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM5 TSMC_10 TSMC_9 VDDI VDDI pch_svt_mac l=20n nfin=4 m=1 
MP10<0> TSMC_12 TSMC_16 TSMC_5 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP10<1> TSMC_12 TSMC_17 TSMC_6 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP10<2> TSMC_12 TSMC_18 TSMC_7 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP10<3> TSMC_12 TSMC_19 TSMC_8 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP3_HDM TSMC_12 TSMC_28 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP22_HDM VDDI TSMC_28 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<0> TSMC_11 TSMC_16 TSMC_1 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<1> TSMC_11 TSMC_17 TSMC_2 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<2> TSMC_11 TSMC_18 TSMC_3 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0<3> TSMC_11 TSMC_19 TSMC_4 VDDI pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_28 TSMC_10 VDDI VDDI pch_svt_mac l=20n nfin=4 m=3 
MM14<0> TSMC_1 TSMC_5 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14<1> TSMC_2 TSMC_6 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14<2> TSMC_3 TSMC_7 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM14<3> TSMC_4 TSMC_8 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<0> TSMC_5 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<1> TSMC_6 TSMC_2 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<2> TSMC_7 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MM13<3> TSMC_8 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
XPRECHARGE<0> TSMC_1 TSMC_5 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW400W20_PRECHARGE_SB_SD 
XPRECHARGE<1> TSMC_2 TSMC_6 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW400W20_PRECHARGE_SB_SD 
XPRECHARGE<2> TSMC_3 TSMC_7 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW400W20_PRECHARGE_SB_SD 
XPRECHARGE<3> TSMC_4 TSMC_8 TSMC_28 VDDI VDDI 
+ S1ALLSVTSW400W20_PRECHARGE_SB_SD 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MIO_M4_SB_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_MIO_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 VSSI TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
XDIN TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_16 TSMC_16 VSSI TSMC_25 TSMC_26 
+ S1ALLSVTSW400W20_DIN_M4_SB_BASE 
XDOUT TSMC_27 TSMC_28 TSMC_29 TSMC_14 TSMC_15 TSMC_16 TSMC_16 VSSI 
+ S1ALLSVTSW400W20_DOUT_SB 
XYPASS TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_27 
+ TSMC_28 TSMC_29 TSMC_13 TSMC_16 VSSI TSMC_25 TSMC_26 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ S1ALLSVTSW400W20_YPASS_M4_SB_NBL_V2 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    CNT_M4_SB_BUF
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_CNT_M4_SB_BUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VSSI 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
XI32 VSSI VSSI TSMC_32 TSMC_4 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=2 n_nfin=10 n_l=20n p_totalM=2 
+ p_nfin=10 p_l=20n 
XI31 VSSI VSSI TSMC_3 TSMC_32 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=10 n_l=20n p_totalM=1 
+ p_nfin=10 p_l=20n 
XWEB_INV VSSI VSSI TSMC_6 TSMC_7 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI29<0> VSSI VSSI TSMC_24 TSMC_28 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI29<1> VSSI VSSI TSMC_25 TSMC_29 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI30 VSSI VSSI TSMC_1 TSMC_2 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
XI28<0> VSSI VSSI TSMC_8 TSMC_16 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<1> VSSI VSSI TSMC_9 TSMC_17 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<2> VSSI VSSI TSMC_10 TSMC_18 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<3> VSSI VSSI TSMC_11 TSMC_19 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<4> VSSI VSSI TSMC_12 TSMC_20 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<5> VSSI VSSI TSMC_13 TSMC_21 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<6> VSSI VSSI TSMC_14 TSMC_22 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI28<7> VSSI VSSI TSMC_15 TSMC_23 TSMC_5 TSMC_5 
+ S1ALLSVTSW400W20_inv_lvt_mac_pcell_6 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    DIODE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_DIODE TSMC_1 TSMC_2 TSMC_3 
MMDIODE TSMC_1 TSMC_2 TSMC_1 TSMC_3 nch_lvt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MCB_D0907_OFFCELL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_MCB_D0907_OFFCELL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
Mpu11 TSMC_9 TSMC_10 TSMC_3 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu21 TSMC_10 TSMC_9 TSMC_8 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_11 TSMC_12 TSMC_3 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu20 TSMC_12 TSMC_11 TSMC_7 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpg21 TSMC_13 TSMC_5 TSMC_10 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd11 TSMC_9 TSMC_10 TSMC_14 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_4 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_12 TSMC_11 TSMC_4 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg11 TSMC_1 TSMC_4 TSMC_9 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_13 TSMC_6 TSMC_12 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_4 TSMC_11 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_11 TSMC_12 TSMC_14 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    LOGIC_D0907_TRKWL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_LOGIC_D0907_TRKWL TSMC_1 TSMC_2 
MM2 TSMC_1 TSMC_2 TSMC_1 TSMC_1 nch_svt_mac l=20n nfin=4 m=1 
MM1 TSMC_1 TSMC_2 TSMC_1 TSMC_1 nch_svt_mac l=20n nfin=4 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MCB_D0907_ONCELL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_MCB_D0907_ONCELL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
Mpd11 TSMC_9 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg21 TSMC_11 TSMC_7 TSMC_10 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_12 TSMC_13 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg11 TSMC_1 TSMC_2 TSMC_9 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_13 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_13 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_11 TSMC_8 TSMC_12 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpu11 TSMC_9 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_13 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: N16FF_SPSB_LEAFCELL
* Cell Name:    MCB_D0907_ONCELL_ISO
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW400W20_MCB_D0907_ONCELL_ISO TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
Mpg11 TSMC_1 TSMC_2 TSMC_10 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd11 TSMC_10 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_11 TSMC_10 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg21 TSMC_12 TSMC_8 TSMC_11 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_13 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_14 TSMC_13 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_13 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_12 TSMC_7 TSMC_14 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpu11 TSMC_10 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_13 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu20 TSMC_15 TSMC_13 TSMC_9 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS




**** End of leaf cells

.SUBCKT S1ALLSVTSW400W20_MCB_ARR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDDAI VDDI VSSI TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 
+ TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 
+ TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 
+ TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 
+ TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
XMCB_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_9 TSMC_10 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_11 TSMC_12 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_13 TSMC_14 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_15 TSMC_16 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI VSSI 
+ TSMC_17 TSMC_18 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_5 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_19 TSMC_20 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_21 TSMC_22 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_7 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_23 TSMC_24 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_25 TSMC_26 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_9 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_27 TSMC_28 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_10 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_29 TSMC_30 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_11 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_31 TSMC_32 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_12 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_33 TSMC_34 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_13 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_35 TSMC_36 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_14 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_37 TSMC_38 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_15 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_39 TSMC_40 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_16 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_41 TSMC_42 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_17 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_43 TSMC_44 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_18 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_45 TSMC_46 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_19 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_47 TSMC_48 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_20 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_49 TSMC_50 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_21 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_51 TSMC_52 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_22 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_53 TSMC_54 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_23 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_55 TSMC_56 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_24 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_57 TSMC_58 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_25 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_59 TSMC_60 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_26 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_61 TSMC_62 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_27 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_63 TSMC_64 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_28 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_65 TSMC_66 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_29 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_67 TSMC_68 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_30 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_69 TSMC_70 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_31 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_71 TSMC_72 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_32 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_73 TSMC_74 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_33 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_75 TSMC_76 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_34 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_77 TSMC_78 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_35 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_79 TSMC_80 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_36 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_81 TSMC_82 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_37 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_83 TSMC_84 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_38 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_85 TSMC_86 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_39 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_87 TSMC_88 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_40 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_89 TSMC_90 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_41 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_91 TSMC_92 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_42 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_93 TSMC_94 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_43 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_95 TSMC_96 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_44 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_97 TSMC_98 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_45 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_99 TSMC_100 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_46 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_101 TSMC_102 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_47 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_103 TSMC_104 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_48 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_105 TSMC_106 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_49 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_107 TSMC_108 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_50 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_109 TSMC_110 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_51 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_111 TSMC_112 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_52 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_113 TSMC_114 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_53 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_115 TSMC_116 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_54 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_117 TSMC_118 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_55 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_119 TSMC_120 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_56 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_121 TSMC_122 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_57 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_123 TSMC_124 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_58 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_125 TSMC_126 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_59 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_127 TSMC_128 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_60 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_129 TSMC_130 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_61 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_131 TSMC_132 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_62 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_133 TSMC_134 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_63 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_135 TSMC_136 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_64 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_137 TSMC_138 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_65 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_139 TSMC_140 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_66 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_141 TSMC_142 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_67 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_143 TSMC_144 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_68 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_145 TSMC_146 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_69 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_147 TSMC_148 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_70 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_149 TSMC_150 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_71 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_151 TSMC_152 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_72 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_153 TSMC_154 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_73 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_155 TSMC_156 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_74 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_157 TSMC_158 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_75 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_159 TSMC_160 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_76 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_161 TSMC_162 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_77 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_163 TSMC_164 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_78 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_165 TSMC_166 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_79 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_167 TSMC_168 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_80 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_169 TSMC_170 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_81 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_171 TSMC_172 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_82 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_173 TSMC_174 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_83 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_175 TSMC_176 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_84 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_177 TSMC_178 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_85 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_179 TSMC_180 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_86 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_181 TSMC_182 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_87 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_183 TSMC_184 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_88 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_185 TSMC_186 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_89 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_187 TSMC_188 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_90 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_189 TSMC_190 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_91 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_191 TSMC_192 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_92 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_193 TSMC_194 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_93 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_195 TSMC_196 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_94 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_197 TSMC_198 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_95 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_199 TSMC_200 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_96 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_201 TSMC_202 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_97 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_203 TSMC_204 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_98 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_205 TSMC_206 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_99 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_207 TSMC_208 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_100 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_209 TSMC_210 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_101 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_211 TSMC_212 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_102 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_213 TSMC_214 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_103 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_215 TSMC_216 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_104 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_217 TSMC_218 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_105 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_219 TSMC_220 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_106 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_221 TSMC_222 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_107 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_223 TSMC_224 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_108 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_225 TSMC_226 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_109 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_227 TSMC_228 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_110 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_229 TSMC_230 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_111 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_231 TSMC_232 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_112 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_233 TSMC_234 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_113 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_235 TSMC_236 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_114 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_237 TSMC_238 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_115 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_239 TSMC_240 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_116 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_241 TSMC_242 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_117 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_243 TSMC_244 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_118 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_245 TSMC_246 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_119 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_247 TSMC_248 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_120 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_249 TSMC_250 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_121 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_251 TSMC_252 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_122 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_253 TSMC_254 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_123 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_255 TSMC_256 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_124 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_257 TSMC_258 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_125 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_259 TSMC_260 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_126 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_261 TSMC_262 S1ALLSVTSW400W20_MCB_2X4_SD 
XMCB_127 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDDAI VDDI 
+ VSSI TSMC_263 TSMC_264 S1ALLSVTSW400W20_MCB_2X4_SD 
.ENDS

.SUBCKT S1ALLSVTSW400W20_TRACKING_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 VDDI VSSI TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 
+ TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 
+ TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 
+ TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 
+ TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 
+ TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 
+ TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 
+ TSMC_322 TSMC_323 
XTKBL_ON_CELL_0 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_321 
+ TSMC_322 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_1 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_319 
+ TSMC_320 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_2 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_317 
+ TSMC_318 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_3 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_315 
+ TSMC_316 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_4 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_313 
+ TSMC_314 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_5 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_311 
+ TSMC_312 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_6 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_309 
+ TSMC_310 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_7 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_307 
+ TSMC_308 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_8 TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_305 
+ TSMC_306 S1ALLSVTSW400W20_MCB_D0907_ONCELL 
XTKBL_ON_CELL_ISO TSMC_65 TSMC_323 TSMC_323 VDDI TSMC_66 VSSI TSMC_303 TSMC_304 
+ TSMC_324 S1ALLSVTSW400W20_MCB_D0907_ONCELL_ISO 
XTKBL_OFF_CELL_10 TSMC_65 VDDI TSMC_66 VSSI TSMC_301 TSMC_302 TSMC_324 
+ TSMC_325 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_11 TSMC_65 VDDI TSMC_66 VSSI TSMC_299 TSMC_300 TSMC_325 
+ TSMC_326 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_12 TSMC_65 VDDI TSMC_66 VSSI TSMC_297 TSMC_298 TSMC_326 
+ TSMC_327 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_13 TSMC_65 VDDI TSMC_66 VSSI TSMC_295 TSMC_296 TSMC_327 
+ TSMC_328 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_14 TSMC_65 VDDI TSMC_66 VSSI TSMC_293 TSMC_294 TSMC_328 
+ TSMC_329 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_15 TSMC_65 VDDI TSMC_66 VSSI TSMC_291 TSMC_292 TSMC_329 
+ TSMC_330 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_16 TSMC_65 VDDI TSMC_66 VSSI TSMC_289 TSMC_290 TSMC_330 
+ TSMC_331 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_17 TSMC_65 VDDI TSMC_66 VSSI TSMC_287 TSMC_288 TSMC_331 
+ TSMC_332 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_18 TSMC_65 VDDI TSMC_66 VSSI TSMC_285 TSMC_286 TSMC_332 
+ TSMC_333 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_19 TSMC_65 VDDI TSMC_66 VSSI TSMC_283 TSMC_284 TSMC_333 
+ TSMC_334 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_20 TSMC_65 VDDI TSMC_66 VSSI TSMC_281 TSMC_282 TSMC_334 
+ TSMC_335 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_21 TSMC_65 VDDI TSMC_66 VSSI TSMC_279 TSMC_280 TSMC_335 
+ TSMC_336 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_22 TSMC_65 VDDI TSMC_66 VSSI TSMC_277 TSMC_278 TSMC_336 
+ TSMC_337 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_23 TSMC_65 VDDI TSMC_66 VSSI TSMC_275 TSMC_276 TSMC_337 
+ TSMC_338 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_24 TSMC_65 VDDI TSMC_66 VSSI TSMC_273 TSMC_274 TSMC_338 
+ TSMC_339 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_25 TSMC_65 VDDI TSMC_66 VSSI TSMC_271 TSMC_272 TSMC_339 
+ TSMC_340 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_26 TSMC_65 VDDI TSMC_66 VSSI TSMC_269 TSMC_270 TSMC_340 
+ TSMC_341 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_27 TSMC_65 VDDI TSMC_66 VSSI TSMC_267 TSMC_268 TSMC_341 
+ TSMC_342 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_28 TSMC_65 VDDI TSMC_66 VSSI TSMC_265 TSMC_266 TSMC_342 
+ TSMC_343 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_29 TSMC_65 VDDI TSMC_66 VSSI TSMC_263 TSMC_264 TSMC_343 
+ TSMC_344 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_30 TSMC_65 VDDI TSMC_66 VSSI TSMC_261 TSMC_262 TSMC_344 
+ TSMC_345 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_31 TSMC_65 VDDI TSMC_66 VSSI TSMC_259 TSMC_260 TSMC_345 
+ TSMC_346 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_32 TSMC_65 VDDI TSMC_66 VSSI TSMC_257 TSMC_258 TSMC_346 
+ TSMC_347 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_33 TSMC_65 VDDI TSMC_66 VSSI TSMC_255 TSMC_256 TSMC_347 
+ TSMC_348 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_34 TSMC_65 VDDI TSMC_66 VSSI TSMC_253 TSMC_254 TSMC_348 
+ TSMC_349 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_35 TSMC_65 VDDI TSMC_66 VSSI TSMC_251 TSMC_252 TSMC_349 
+ TSMC_350 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_36 TSMC_65 VDDI TSMC_66 VSSI TSMC_249 TSMC_250 TSMC_350 
+ TSMC_351 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_37 TSMC_65 VDDI TSMC_66 VSSI TSMC_247 TSMC_248 TSMC_351 
+ TSMC_352 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_38 TSMC_65 VDDI TSMC_66 VSSI TSMC_245 TSMC_246 TSMC_352 
+ TSMC_353 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_39 TSMC_65 VDDI TSMC_66 VSSI TSMC_243 TSMC_244 TSMC_353 
+ TSMC_354 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_40 TSMC_65 VDDI TSMC_66 VSSI TSMC_241 TSMC_242 TSMC_354 
+ TSMC_355 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_41 TSMC_65 VDDI TSMC_66 VSSI TSMC_239 TSMC_240 TSMC_355 
+ TSMC_356 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_42 TSMC_65 VDDI TSMC_66 VSSI TSMC_237 TSMC_238 TSMC_356 
+ TSMC_357 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_43 TSMC_65 VDDI TSMC_66 VSSI TSMC_235 TSMC_236 TSMC_357 
+ TSMC_358 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_44 TSMC_65 VDDI TSMC_66 VSSI TSMC_233 TSMC_234 TSMC_358 
+ TSMC_359 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_45 TSMC_65 VDDI TSMC_66 VSSI TSMC_231 TSMC_232 TSMC_359 
+ TSMC_360 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_46 TSMC_65 VDDI TSMC_66 VSSI TSMC_229 TSMC_230 TSMC_360 
+ TSMC_361 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_47 TSMC_65 VDDI TSMC_66 VSSI TSMC_227 TSMC_228 TSMC_361 
+ TSMC_362 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_48 TSMC_65 VDDI TSMC_66 VSSI TSMC_225 TSMC_226 TSMC_362 
+ TSMC_363 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_49 TSMC_65 VDDI TSMC_66 VSSI TSMC_223 TSMC_224 TSMC_363 
+ TSMC_364 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_50 TSMC_65 VDDI TSMC_66 VSSI TSMC_221 TSMC_222 TSMC_364 
+ TSMC_365 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_51 TSMC_65 VDDI TSMC_66 VSSI TSMC_219 TSMC_220 TSMC_365 
+ TSMC_366 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_52 TSMC_65 VDDI TSMC_66 VSSI TSMC_217 TSMC_218 TSMC_366 
+ TSMC_367 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_53 TSMC_65 VDDI TSMC_66 VSSI TSMC_215 TSMC_216 TSMC_367 
+ TSMC_368 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_54 TSMC_65 VDDI TSMC_66 VSSI TSMC_213 TSMC_214 TSMC_368 
+ TSMC_369 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_55 TSMC_65 VDDI TSMC_66 VSSI TSMC_211 TSMC_212 TSMC_369 
+ TSMC_370 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_56 TSMC_65 VDDI TSMC_66 VSSI TSMC_209 TSMC_210 TSMC_370 
+ TSMC_371 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_57 TSMC_65 VDDI TSMC_66 VSSI TSMC_207 TSMC_208 TSMC_371 
+ TSMC_372 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_58 TSMC_65 VDDI TSMC_66 VSSI TSMC_205 TSMC_206 TSMC_372 
+ TSMC_373 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_59 TSMC_65 VDDI TSMC_66 VSSI TSMC_203 TSMC_204 TSMC_373 
+ TSMC_374 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_60 TSMC_65 VDDI TSMC_66 VSSI TSMC_201 TSMC_202 TSMC_374 
+ TSMC_375 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_61 TSMC_65 VDDI TSMC_66 VSSI TSMC_199 TSMC_200 TSMC_375 
+ TSMC_376 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_62 TSMC_65 VDDI TSMC_66 VSSI TSMC_197 TSMC_198 TSMC_376 
+ TSMC_377 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_63 TSMC_65 VDDI TSMC_66 VSSI TSMC_195 TSMC_196 TSMC_377 
+ TSMC_378 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_64 TSMC_65 VDDI TSMC_66 VSSI TSMC_193 TSMC_194 TSMC_378 
+ TSMC_379 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_65 TSMC_65 VDDI TSMC_66 VSSI TSMC_191 TSMC_192 TSMC_379 
+ TSMC_380 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_66 TSMC_65 VDDI TSMC_66 VSSI TSMC_189 TSMC_190 TSMC_380 
+ TSMC_381 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_67 TSMC_65 VDDI TSMC_66 VSSI TSMC_187 TSMC_188 TSMC_381 
+ TSMC_382 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_68 TSMC_65 VDDI TSMC_66 VSSI TSMC_185 TSMC_186 TSMC_382 
+ TSMC_383 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_69 TSMC_65 VDDI TSMC_66 VSSI TSMC_183 TSMC_184 TSMC_383 
+ TSMC_384 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_70 TSMC_65 VDDI TSMC_66 VSSI TSMC_181 TSMC_182 TSMC_384 
+ TSMC_385 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_71 TSMC_65 VDDI TSMC_66 VSSI TSMC_179 TSMC_180 TSMC_385 
+ TSMC_386 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_72 TSMC_65 VDDI TSMC_66 VSSI TSMC_177 TSMC_178 TSMC_386 
+ TSMC_387 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_73 TSMC_65 VDDI TSMC_66 VSSI TSMC_175 TSMC_176 TSMC_387 
+ TSMC_388 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_74 TSMC_65 VDDI TSMC_66 VSSI TSMC_173 TSMC_174 TSMC_388 
+ TSMC_389 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_75 TSMC_65 VDDI TSMC_66 VSSI TSMC_171 TSMC_172 TSMC_389 
+ TSMC_390 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_76 TSMC_65 VDDI TSMC_66 VSSI TSMC_169 TSMC_170 TSMC_390 
+ TSMC_391 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_77 TSMC_65 VDDI TSMC_66 VSSI TSMC_167 TSMC_168 TSMC_391 
+ TSMC_392 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_78 TSMC_65 VDDI TSMC_66 VSSI TSMC_165 TSMC_166 TSMC_392 
+ TSMC_393 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_79 TSMC_65 VDDI TSMC_66 VSSI TSMC_163 TSMC_164 TSMC_393 
+ TSMC_394 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_80 TSMC_65 VDDI TSMC_66 VSSI TSMC_161 TSMC_162 TSMC_394 
+ TSMC_395 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_81 TSMC_65 VDDI TSMC_66 VSSI TSMC_159 TSMC_160 TSMC_395 
+ TSMC_396 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_82 TSMC_65 VDDI TSMC_66 VSSI TSMC_157 TSMC_158 TSMC_396 
+ TSMC_397 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_83 TSMC_65 VDDI TSMC_66 VSSI TSMC_155 TSMC_156 TSMC_397 
+ TSMC_398 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_84 TSMC_65 VDDI TSMC_66 VSSI TSMC_153 TSMC_154 TSMC_398 
+ TSMC_399 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_85 TSMC_65 VDDI TSMC_66 VSSI TSMC_151 TSMC_152 TSMC_399 
+ TSMC_400 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_86 TSMC_65 VDDI TSMC_66 VSSI TSMC_149 TSMC_150 TSMC_400 
+ TSMC_401 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_87 TSMC_65 VDDI TSMC_66 VSSI TSMC_147 TSMC_148 TSMC_401 
+ TSMC_402 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_88 TSMC_65 VDDI TSMC_66 VSSI TSMC_145 TSMC_146 TSMC_402 
+ TSMC_403 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_89 TSMC_65 VDDI TSMC_66 VSSI TSMC_143 TSMC_144 TSMC_403 
+ TSMC_404 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_90 TSMC_65 VDDI TSMC_66 VSSI TSMC_141 TSMC_142 TSMC_404 
+ TSMC_405 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_91 TSMC_65 VDDI TSMC_66 VSSI TSMC_139 TSMC_140 TSMC_405 
+ TSMC_406 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_92 TSMC_65 VDDI TSMC_66 VSSI TSMC_137 TSMC_138 TSMC_406 
+ TSMC_407 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_93 TSMC_65 VDDI TSMC_66 VSSI TSMC_135 TSMC_136 TSMC_407 
+ TSMC_408 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_94 TSMC_65 VDDI TSMC_66 VSSI TSMC_133 TSMC_134 TSMC_408 
+ TSMC_409 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_95 TSMC_65 VDDI TSMC_66 VSSI TSMC_131 TSMC_132 TSMC_409 
+ TSMC_410 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_96 TSMC_65 VDDI TSMC_66 VSSI TSMC_129 TSMC_130 TSMC_410 
+ TSMC_411 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_97 TSMC_65 VDDI TSMC_66 VSSI TSMC_127 TSMC_128 TSMC_411 
+ TSMC_412 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_98 TSMC_65 VDDI TSMC_66 VSSI TSMC_125 TSMC_126 TSMC_412 
+ TSMC_413 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_99 TSMC_65 VDDI TSMC_66 VSSI TSMC_123 TSMC_124 TSMC_413 
+ TSMC_414 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_100 TSMC_65 VDDI TSMC_66 VSSI TSMC_121 TSMC_122 
+ TSMC_414 TSMC_415 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_101 TSMC_65 VDDI TSMC_66 VSSI TSMC_119 TSMC_120 
+ TSMC_415 TSMC_416 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_102 TSMC_65 VDDI TSMC_66 VSSI TSMC_117 TSMC_118 
+ TSMC_416 TSMC_417 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_103 TSMC_65 VDDI TSMC_66 VSSI TSMC_115 TSMC_116 
+ TSMC_417 TSMC_418 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_104 TSMC_65 VDDI TSMC_66 VSSI TSMC_113 TSMC_114 
+ TSMC_418 TSMC_419 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_105 TSMC_65 VDDI TSMC_66 VSSI TSMC_111 TSMC_112 
+ TSMC_419 TSMC_420 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_106 TSMC_65 VDDI TSMC_66 VSSI TSMC_109 TSMC_110 
+ TSMC_420 TSMC_421 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_107 TSMC_65 VDDI TSMC_66 VSSI TSMC_107 TSMC_108 
+ TSMC_421 TSMC_422 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_108 TSMC_65 VDDI TSMC_66 VSSI TSMC_105 TSMC_106 
+ TSMC_422 TSMC_423 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_109 TSMC_65 VDDI TSMC_66 VSSI TSMC_103 TSMC_104 
+ TSMC_423 TSMC_424 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_110 TSMC_65 VDDI TSMC_66 VSSI TSMC_101 TSMC_102 
+ TSMC_424 TSMC_425 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_111 TSMC_65 VDDI TSMC_66 VSSI TSMC_99 TSMC_100 TSMC_425 
+ TSMC_426 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_112 TSMC_65 VDDI TSMC_66 VSSI TSMC_97 TSMC_98 TSMC_426 
+ TSMC_427 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_113 TSMC_65 VDDI TSMC_66 VSSI TSMC_95 TSMC_96 TSMC_427 
+ TSMC_428 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_114 TSMC_65 VDDI TSMC_66 VSSI TSMC_93 TSMC_94 TSMC_428 
+ TSMC_429 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_115 TSMC_65 VDDI TSMC_66 VSSI TSMC_91 TSMC_92 TSMC_429 
+ TSMC_430 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_116 TSMC_65 VDDI TSMC_66 VSSI TSMC_89 TSMC_90 TSMC_430 
+ TSMC_431 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_117 TSMC_65 VDDI TSMC_66 VSSI TSMC_87 TSMC_88 TSMC_431 
+ TSMC_432 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_118 TSMC_65 VDDI TSMC_66 VSSI TSMC_85 TSMC_86 TSMC_432 
+ TSMC_433 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_119 TSMC_65 VDDI TSMC_66 VSSI TSMC_83 TSMC_84 TSMC_433 
+ TSMC_434 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_120 TSMC_65 VDDI TSMC_66 VSSI TSMC_81 TSMC_82 TSMC_434 
+ TSMC_435 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_121 TSMC_65 VDDI TSMC_66 VSSI TSMC_79 TSMC_80 TSMC_435 
+ TSMC_436 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_122 TSMC_65 VDDI TSMC_66 VSSI TSMC_77 TSMC_78 TSMC_436 
+ TSMC_437 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_123 TSMC_65 VDDI TSMC_66 VSSI TSMC_75 TSMC_76 TSMC_437 
+ TSMC_438 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_124 TSMC_65 VDDI TSMC_66 VSSI TSMC_73 TSMC_74 TSMC_438 
+ TSMC_439 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_125 TSMC_65 VDDI TSMC_66 VSSI TSMC_71 TSMC_72 TSMC_439 
+ TSMC_440 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_126 TSMC_65 VDDI TSMC_66 VSSI TSMC_69 TSMC_70 TSMC_440 
+ TSMC_441 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTKBL_OFF_CELL_127 TSMC_65 VDDI TSMC_66 VSSI TSMC_67 TSMC_68 TSMC_441 
+ TSMC_442 S1ALLSVTSW400W20_MCB_D0907_OFFCELL 
XTRKWL_CELL_0 VSSI TSMC_323 S1ALLSVTSW400W20_LOGIC_D0907_TRKWL 
XTRKWL_CELL_1 VSSI TSMC_323 S1ALLSVTSW400W20_LOGIC_D0907_TRKWL 
XTRKWL_CELL_2 VSSI TSMC_323 S1ALLSVTSW400W20_LOGIC_D0907_TRKWL 
.ENDS

.SUBCKT S1ALLSVTSW400W20_MIO_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 VSSI 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
XMIO_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_24 TSMC_11 TSMC_25 VSSI TSMC_13 TSMC_14 TSMC_15 VSSI TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ S1ALLSVTSW400W20_MIO_M4_SB_BASE 
XMIO_MX_SB_BUF TSMC_10 TSMC_24 TSMC_12 TSMC_25 TSMC_15 VSSI 
+ S1ALLSVTSW400W20_MIO_M4_SB_BUF 
.ENDS

.SUBCKT S1ALLSVTSW400W20_CNT_M4_SB TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 VSSI TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
XCNT_M4_SB_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_62 TSMC_5 TSMC_6 TSMC_63 TSMC_7 
+ TSMC_64 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 VSSI TSMC_65 
+ TSMC_66 TSMC_47 TSMC_48 TSMC_49 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ S1ALLSVTSW400W20_CNT_M4_SB_BASE 
XCNT_MX_SB_BUF TSMC_4 TSMC_62 TSMC_7 TSMC_64 TSMC_45 VSSI TSMC_46 TSMC_65 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_58 
+ TSMC_59 TSMC_60 TSMC_61 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ S1ALLSVTSW400W20_CNT_M4_SB_BUF 
.ENDS

.SUBCKT TS1N16FFCLLSVTA1024X32M4SW D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] D[8] 
+ D[9] D[10] D[11] D[12] D[13] D[14] D[15] D[16] D[17] D[18] D[19] D[20] D[21] 
+ D[22] D[23] D[24] D[25] D[26] D[27] D[28] D[29] D[30] D[31] BWEB[0] BWEB[1] 
+ BWEB[2] BWEB[3] BWEB[4] BWEB[5] BWEB[6] BWEB[7] BWEB[8] BWEB[9] BWEB[10] 
+ BWEB[11] BWEB[12] BWEB[13] BWEB[14] BWEB[15] BWEB[16] BWEB[17] BWEB[18] 
+ BWEB[19] BWEB[20] BWEB[21] BWEB[22] BWEB[23] BWEB[24] BWEB[25] BWEB[26] 
+ BWEB[27] BWEB[28] BWEB[29] BWEB[30] BWEB[31] A[0] A[1] A[2] A[3] A[4] A[5] 
+ A[6] A[7] A[8] A[9] Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] 
+ Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18] Q[19] Q[20] Q[21] Q[22] Q[23] 
+ Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] CEB CLK WEB RTSEL[1] RTSEL[0] 
+ WTSEL[1] WTSEL[0] VDD VSS 
XMCB256X4_L_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDD VDD 
+ VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 
+ TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 
+ TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 
+ TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 
+ TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 
+ TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 
+ TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 
+ TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 
+ TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 
+ TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 
+ TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 
+ TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 
+ TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 
+ TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 
+ TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_1 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_2 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 
+ TSMC_280 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_3 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 
+ TSMC_288 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_4 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 
+ TSMC_296 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_5 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_6 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
+ TSMC_312 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_7 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_8 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 
+ TSMC_328 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_9 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 
+ TSMC_336 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_10 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 
+ TSMC_344 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_11 TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 
+ TSMC_352 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_12 TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 
+ TSMC_360 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_13 TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_14 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_L_15 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 
+ TSMC_384 VDD VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 
+ TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 
+ TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 
+ TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_16 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 
+ TSMC_392 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_17 TSMC_649 TSMC_650 TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 
+ TSMC_656 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_18 TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 TSMC_663 
+ TSMC_664 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_19 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 TSMC_671 
+ TSMC_672 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_20 TSMC_673 TSMC_674 TSMC_675 TSMC_676 TSMC_677 TSMC_678 TSMC_679 
+ TSMC_680 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_21 TSMC_681 TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 TSMC_687 
+ TSMC_688 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_22 TSMC_689 TSMC_690 TSMC_691 TSMC_692 TSMC_693 TSMC_694 TSMC_695 
+ TSMC_696 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_23 TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_701 TSMC_702 TSMC_703 
+ TSMC_704 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_24 TSMC_705 TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 TSMC_711 
+ TSMC_712 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_25 TSMC_713 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 
+ TSMC_719 TSMC_720 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_26 TSMC_721 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_727 TSMC_728 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_27 TSMC_729 TSMC_730 TSMC_731 TSMC_732 TSMC_733 TSMC_734 
+ TSMC_735 TSMC_736 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_28 TSMC_737 TSMC_738 TSMC_739 TSMC_740 TSMC_741 TSMC_742 
+ TSMC_743 TSMC_744 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_29 TSMC_745 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 
+ TSMC_751 TSMC_752 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_30 TSMC_753 TSMC_754 TSMC_755 TSMC_756 TSMC_757 TSMC_758 
+ TSMC_759 TSMC_760 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XMCB256X4_R_31 TSMC_761 TSMC_762 TSMC_763 TSMC_764 TSMC_765 TSMC_766 
+ TSMC_767 TSMC_768 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 
+ TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 
+ TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 
+ TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 
+ TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 
+ S1ALLSVTSW400W20_MCB_ARR 
XXDRV_STRAP_BT_SB_0 TSMC_769 TSMC_770 VDD VSS 
+ S1ALLSVTSW400W20_XDRV_STRAP_BT_SB 
XXDRV_LA512_SB_0 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_775 TSMC_776 
+ TSMC_777 TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_782 TSMC_783 
+ TSMC_784 TSMC_785 TSMC_786 TSMC_787 TSMC_788 TSMC_789 VDD VSS 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_1 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_794 TSMC_795 
+ TSMC_796 TSMC_797 TSMC_779 TSMC_798 TSMC_799 TSMC_800 TSMC_801 
+ TSMC_802 TSMC_803 TSMC_804 TSMC_805 TSMC_806 TSMC_807 VDD VSS 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_2 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_808 TSMC_809 
+ TSMC_810 TSMC_811 TSMC_812 TSMC_813 TSMC_814 TSMC_815 TSMC_816 
+ TSMC_817 TSMC_818 TSMC_819 TSMC_820 TSMC_821 TSMC_822 VDD VSS 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_401 TSMC_402 TSMC_403 TSMC_404 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_3 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_823 TSMC_824 
+ TSMC_825 TSMC_826 TSMC_812 TSMC_827 TSMC_828 TSMC_829 TSMC_830 
+ TSMC_831 TSMC_832 TSMC_833 TSMC_834 TSMC_835 TSMC_836 VDD VSS 
+ TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_405 TSMC_406 TSMC_407 TSMC_408 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_4 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_837 TSMC_838 
+ TSMC_839 TSMC_840 TSMC_841 TSMC_842 TSMC_843 TSMC_844 TSMC_845 
+ TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 VDD VSS 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_409 TSMC_410 TSMC_411 TSMC_412 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_5 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_852 TSMC_853 
+ TSMC_854 TSMC_855 TSMC_841 TSMC_856 TSMC_857 TSMC_858 TSMC_859 
+ TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 VDD VSS 
+ TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_413 TSMC_414 TSMC_415 TSMC_416 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_6 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_866 TSMC_867 
+ TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 TSMC_873 TSMC_874 
+ TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 TSMC_880 VDD VSS 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_417 TSMC_418 TSMC_419 TSMC_420 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_7 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_881 TSMC_882 
+ TSMC_883 TSMC_884 TSMC_870 TSMC_885 TSMC_886 TSMC_887 TSMC_888 
+ TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 VDD VSS 
+ TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_421 TSMC_422 TSMC_423 TSMC_424 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_8 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_895 TSMC_896 
+ TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 TSMC_902 TSMC_903 
+ TSMC_904 TSMC_905 TSMC_906 TSMC_907 TSMC_908 TSMC_909 VDD VSS 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_425 TSMC_426 TSMC_427 TSMC_428 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_9 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_910 TSMC_911 
+ TSMC_912 TSMC_913 TSMC_899 TSMC_914 TSMC_915 TSMC_916 TSMC_917 
+ TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 TSMC_923 VDD VSS 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_769 TSMC_770 S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_10 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_924 
+ TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 TSMC_930 TSMC_931 
+ TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 TSMC_937 
+ TSMC_938 VDD VSS TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_433 TSMC_434 
+ TSMC_435 TSMC_436 TSMC_769 TSMC_770 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_11 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_939 
+ TSMC_940 TSMC_941 TSMC_942 TSMC_928 TSMC_943 TSMC_944 TSMC_945 
+ TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 TSMC_951 
+ TSMC_952 VDD VSS TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_437 TSMC_438 
+ TSMC_439 TSMC_440 TSMC_769 TSMC_770 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_12 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_953 
+ TSMC_954 TSMC_955 TSMC_956 TSMC_957 TSMC_958 TSMC_959 TSMC_960 
+ TSMC_961 TSMC_962 TSMC_963 TSMC_964 TSMC_965 TSMC_966 
+ TSMC_967 VDD VSS TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_441 TSMC_442 
+ TSMC_443 TSMC_444 TSMC_769 TSMC_770 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_13 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_968 
+ TSMC_969 TSMC_970 TSMC_971 TSMC_957 TSMC_972 TSMC_973 TSMC_974 
+ TSMC_975 TSMC_976 TSMC_977 TSMC_978 TSMC_979 TSMC_980 
+ TSMC_981 VDD VSS TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_445 TSMC_446 
+ TSMC_447 TSMC_448 TSMC_769 TSMC_770 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_14 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_982 
+ TSMC_983 TSMC_984 TSMC_985 TSMC_986 TSMC_987 TSMC_988 TSMC_989 
+ TSMC_990 TSMC_991 TSMC_992 TSMC_993 TSMC_994 TSMC_995 
+ TSMC_996 VDD VSS TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_449 TSMC_450 
+ TSMC_451 TSMC_452 TSMC_769 TSMC_770 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_15 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_997 
+ TSMC_998 TSMC_999 TSMC_1000 TSMC_986 TSMC_1001 TSMC_1002 TSMC_1003 
+ TSMC_1004 TSMC_1005 TSMC_1006 TSMC_1007 TSMC_1008 
+ TSMC_1009 TSMC_1010 VDD VSS TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_453 
+ TSMC_454 TSMC_455 TSMC_456 TSMC_769 TSMC_770 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_STRAP_SB_16 TSMC_1011 TSMC_1012 VDD VSS 
+ S1ALLSVTSW400W20_XDRV_STRAP_SB 
XXDRV_LA512_SB_16 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1013 
+ TSMC_1014 TSMC_1015 TSMC_1016 TSMC_779 TSMC_1017 TSMC_1018 
+ TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 
+ TSMC_1025 TSMC_1026 VDD VSS TSMC_73 TSMC_74 TSMC_75 TSMC_76 
+ TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_17 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1027 
+ TSMC_1028 TSMC_1029 TSMC_1030 TSMC_779 TSMC_1031 TSMC_1032 
+ TSMC_1033 TSMC_1034 TSMC_1035 TSMC_1036 TSMC_1037 TSMC_1038 
+ TSMC_1039 TSMC_1040 VDD VSS TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_18 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1041 
+ TSMC_1042 TSMC_1043 TSMC_1044 TSMC_812 TSMC_1045 TSMC_1046 
+ TSMC_1047 TSMC_1048 TSMC_1049 TSMC_1050 TSMC_1051 TSMC_1052 
+ TSMC_1053 TSMC_1054 VDD VSS TSMC_81 TSMC_82 TSMC_83 TSMC_84 
+ TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_19 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_812 TSMC_1059 TSMC_1060 
+ TSMC_1061 TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 
+ TSMC_1067 TSMC_1068 VDD VSS TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_20 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1069 
+ TSMC_1070 TSMC_1071 TSMC_1072 TSMC_841 TSMC_1073 TSMC_1074 
+ TSMC_1075 TSMC_1076 TSMC_1077 TSMC_1078 TSMC_1079 TSMC_1080 
+ TSMC_1081 TSMC_1082 VDD VSS TSMC_89 TSMC_90 TSMC_91 TSMC_92 
+ TSMC_473 TSMC_474 TSMC_475 TSMC_476 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_21 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1083 
+ TSMC_1084 TSMC_1085 TSMC_1086 TSMC_841 TSMC_1087 TSMC_1088 
+ TSMC_1089 TSMC_1090 TSMC_1091 TSMC_1092 TSMC_1093 TSMC_1094 
+ TSMC_1095 TSMC_1096 VDD VSS TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_22 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1097 
+ TSMC_1098 TSMC_1099 TSMC_1100 TSMC_870 TSMC_1101 TSMC_1102 
+ TSMC_1103 TSMC_1104 TSMC_1105 TSMC_1106 TSMC_1107 TSMC_1108 
+ TSMC_1109 TSMC_1110 VDD VSS TSMC_97 TSMC_98 TSMC_99 TSMC_100 
+ TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_23 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1111 
+ TSMC_1112 TSMC_1113 TSMC_1114 TSMC_870 TSMC_1115 TSMC_1116 
+ TSMC_1117 TSMC_1118 TSMC_1119 TSMC_1120 TSMC_1121 TSMC_1122 
+ TSMC_1123 TSMC_1124 VDD VSS TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_24 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1125 
+ TSMC_1126 TSMC_1127 TSMC_1128 TSMC_899 TSMC_1129 TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 TSMC_1138 VDD VSS TSMC_105 TSMC_106 TSMC_107 TSMC_108 
+ TSMC_489 TSMC_490 TSMC_491 TSMC_492 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_25 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1139 
+ TSMC_1140 TSMC_1141 TSMC_1142 TSMC_899 TSMC_1143 TSMC_1144 
+ TSMC_1145 TSMC_1146 TSMC_1147 TSMC_1148 TSMC_1149 TSMC_1150 
+ TSMC_1151 TSMC_1152 VDD VSS TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_26 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1153 
+ TSMC_1154 TSMC_1155 TSMC_1156 TSMC_928 TSMC_1157 TSMC_1158 
+ TSMC_1159 TSMC_1160 TSMC_1161 TSMC_1162 TSMC_1163 TSMC_1164 
+ TSMC_1165 TSMC_1166 VDD VSS TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_27 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1167 
+ TSMC_1168 TSMC_1169 TSMC_1170 TSMC_928 TSMC_1171 TSMC_1172 
+ TSMC_1173 TSMC_1174 TSMC_1175 TSMC_1176 TSMC_1177 TSMC_1178 
+ TSMC_1179 TSMC_1180 VDD VSS TSMC_117 TSMC_118 TSMC_119 TSMC_120 
+ TSMC_501 TSMC_502 TSMC_503 TSMC_504 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_28 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1181 
+ TSMC_1182 TSMC_1183 TSMC_1184 TSMC_957 TSMC_1185 TSMC_1186 
+ TSMC_1187 TSMC_1188 TSMC_1189 TSMC_1190 TSMC_1191 TSMC_1192 
+ TSMC_1193 TSMC_1194 VDD VSS TSMC_121 TSMC_122 TSMC_123 TSMC_124 
+ TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_29 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1195 
+ TSMC_1196 TSMC_1197 TSMC_1198 TSMC_957 TSMC_1199 TSMC_1200 
+ TSMC_1201 TSMC_1202 TSMC_1203 TSMC_1204 TSMC_1205 TSMC_1206 
+ TSMC_1207 TSMC_1208 VDD VSS TSMC_125 TSMC_126 TSMC_127 TSMC_128 
+ TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_30 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1209 
+ TSMC_1210 TSMC_1211 TSMC_1212 TSMC_986 TSMC_1213 TSMC_1214 
+ TSMC_1215 TSMC_1216 TSMC_1217 TSMC_1218 TSMC_1219 TSMC_1220 
+ TSMC_1221 TSMC_1222 VDD VSS TSMC_129 TSMC_130 TSMC_131 TSMC_132 
+ TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_31 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1223 
+ TSMC_1224 TSMC_1225 TSMC_1226 TSMC_986 TSMC_1227 TSMC_1228 
+ TSMC_1229 TSMC_1230 TSMC_1231 TSMC_1232 TSMC_1233 TSMC_1234 
+ TSMC_1235 TSMC_1236 VDD VSS TSMC_133 TSMC_134 TSMC_135 TSMC_136 
+ TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_1011 TSMC_1012 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_STRAP_SB_32 TSMC_1237 TSMC_1238 VDD VSS 
+ S1ALLSVTSW400W20_XDRV_STRAP_SB 
XXDRV_LA512_SB_32 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1239 
+ TSMC_1240 TSMC_1241 TSMC_1242 TSMC_779 TSMC_1243 TSMC_1244 
+ TSMC_1245 TSMC_1246 TSMC_1247 TSMC_1248 TSMC_1249 TSMC_1250 
+ TSMC_1251 TSMC_1252 VDD VSS TSMC_137 TSMC_138 TSMC_139 TSMC_140 
+ TSMC_521 TSMC_522 TSMC_523 TSMC_524 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_33 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_779 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 
+ TSMC_1265 TSMC_1266 VDD VSS TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_34 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_812 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 VDD VSS TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_35 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_812 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 VDD VSS TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_36 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1295 
+ TSMC_1296 TSMC_1297 TSMC_1298 TSMC_841 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 VDD VSS TSMC_153 TSMC_154 TSMC_155 TSMC_156 
+ TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_37 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1309 
+ TSMC_1310 TSMC_1311 TSMC_1312 TSMC_841 TSMC_1313 TSMC_1314 
+ TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 
+ TSMC_1321 TSMC_1322 VDD VSS TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_38 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_870 TSMC_1327 TSMC_1328 
+ TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 
+ TSMC_1335 TSMC_1336 VDD VSS TSMC_161 TSMC_162 TSMC_163 TSMC_164 
+ TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_39 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_870 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 VDD VSS TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_40 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_899 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 VDD VSS TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_41 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1365 
+ TSMC_1366 TSMC_1367 TSMC_1368 TSMC_899 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 VDD VSS TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_557 TSMC_558 TSMC_559 TSMC_560 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_42 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1379 
+ TSMC_1380 TSMC_1381 TSMC_1382 TSMC_928 TSMC_1383 TSMC_1384 
+ TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 
+ TSMC_1391 TSMC_1392 VDD VSS TSMC_177 TSMC_178 TSMC_179 TSMC_180 
+ TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_43 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_928 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 
+ TSMC_1405 TSMC_1406 VDD VSS TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_565 TSMC_566 TSMC_567 TSMC_568 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_44 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_957 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 VDD VSS TSMC_185 TSMC_186 TSMC_187 TSMC_188 
+ TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_45 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_957 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 VDD VSS TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_573 TSMC_574 TSMC_575 TSMC_576 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_46 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1435 
+ TSMC_1436 TSMC_1437 TSMC_1438 TSMC_986 TSMC_1439 TSMC_1440 
+ TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 VDD VSS TSMC_193 TSMC_194 TSMC_195 TSMC_196 
+ TSMC_577 TSMC_578 TSMC_579 TSMC_580 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_47 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_986 TSMC_1453 TSMC_1454 
+ TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 
+ TSMC_1461 TSMC_1462 VDD VSS TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_1237 TSMC_1238 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_STRAP_SB_48 TSMC_1463 TSMC_1464 VDD VSS 
+ S1ALLSVTSW400W20_XDRV_STRAP_SB 
XXDRV_LA512_SB_48 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_779 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 VDD VSS TSMC_201 TSMC_202 TSMC_203 TSMC_204 
+ TSMC_585 TSMC_586 TSMC_587 TSMC_588 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_49 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1479 
+ TSMC_1480 TSMC_1481 TSMC_1482 TSMC_779 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 VDD VSS TSMC_205 TSMC_206 TSMC_207 TSMC_208 
+ TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_50 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_812 TSMC_1497 TSMC_1498 
+ TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ TSMC_1505 TSMC_1506 VDD VSS TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_51 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1507 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_812 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 VDD VSS TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_52 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1521 
+ TSMC_1522 TSMC_1523 TSMC_1524 TSMC_841 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 
+ TSMC_1533 TSMC_1534 VDD VSS TSMC_217 TSMC_218 TSMC_219 TSMC_220 
+ TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_53 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1535 
+ TSMC_1536 TSMC_1537 TSMC_1538 TSMC_841 TSMC_1539 TSMC_1540 
+ TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 TSMC_1546 
+ TSMC_1547 TSMC_1548 VDD VSS TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_605 TSMC_606 TSMC_607 TSMC_608 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_54 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_870 TSMC_1553 TSMC_1554 
+ TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 
+ TSMC_1561 TSMC_1562 VDD VSS TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_55 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_870 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 
+ TSMC_1575 TSMC_1576 VDD VSS TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_56 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_899 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 VDD VSS TSMC_233 TSMC_234 TSMC_235 TSMC_236 
+ TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_57 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1591 
+ TSMC_1592 TSMC_1593 TSMC_1594 TSMC_899 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 VDD VSS TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_621 TSMC_622 TSMC_623 TSMC_624 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_58 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1605 
+ TSMC_1606 TSMC_1607 TSMC_1608 TSMC_928 TSMC_1609 TSMC_1610 
+ TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 
+ TSMC_1617 TSMC_1618 VDD VSS TSMC_241 TSMC_242 TSMC_243 TSMC_244 
+ TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_59 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_928 TSMC_1623 TSMC_1624 
+ TSMC_1625 TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 
+ TSMC_1631 TSMC_1632 VDD VSS TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_629 TSMC_630 TSMC_631 TSMC_632 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_60 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_957 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 VDD VSS TSMC_249 TSMC_250 TSMC_251 TSMC_252 
+ TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_61 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1647 
+ TSMC_1648 TSMC_1649 TSMC_1650 TSMC_957 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 VDD VSS TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_62 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_1661 
+ TSMC_1662 TSMC_1663 TSMC_1664 TSMC_986 TSMC_1665 TSMC_1666 
+ TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 TSMC_1672 
+ TSMC_1673 TSMC_1674 VDD VSS TSMC_257 TSMC_258 TSMC_259 TSMC_260 
+ TSMC_641 TSMC_642 TSMC_643 TSMC_644 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XXDRV_LA512_SB_63 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_986 TSMC_1679 TSMC_1680 
+ TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 
+ TSMC_1687 TSMC_1688 VDD VSS TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_1463 TSMC_1464 
+ S1ALLSVTSW400W20_XDRV_LA512_884_SB 
XTRACKING_XB256X4 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_665 
+ TSMC_666 TSMC_667 TSMC_668 TSMC_673 TSMC_674 TSMC_675 TSMC_676 
+ TSMC_681 TSMC_682 TSMC_683 TSMC_684 TSMC_689 TSMC_690 TSMC_691 
+ TSMC_692 TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_705 TSMC_706 
+ TSMC_707 TSMC_708 TSMC_713 TSMC_714 TSMC_715 TSMC_716 TSMC_721 TSMC_722 
+ TSMC_723 TSMC_724 TSMC_729 TSMC_730 TSMC_731 TSMC_732 TSMC_737 
+ TSMC_738 TSMC_739 TSMC_740 TSMC_745 TSMC_746 TSMC_747 TSMC_748 
+ TSMC_753 TSMC_754 TSMC_755 TSMC_756 TSMC_761 TSMC_762 TSMC_763 
+ TSMC_764 TSMC_1689 VDD VDD VSS TSMC_393 TSMC_394 TSMC_395 TSMC_396 
+ TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 
+ TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 
+ TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 
+ TSMC_447 TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 
+ TSMC_454 TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 TSMC_460 
+ TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 
+ TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 
+ TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 
+ TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 
+ TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 TSMC_524 
+ TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 TSMC_531 
+ TSMC_532 TSMC_533 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 
+ TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 
+ TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 
+ TSMC_553 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 
+ TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 
+ TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_598 TSMC_599 TSMC_600 TSMC_601 
+ TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 
+ TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 
+ TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 
+ TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_1690 
+ S1ALLSVTSW400W20_TRACKING_SB 
XMIOM4_L_0 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_1691 
+ BWEB[0] TSMC_1692 D[0] Q[0] TSMC_1693 VDD VSS TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_1 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_265 TSMC_266 TSMC_267 
+ TSMC_268 TSMC_1691 BWEB[1] TSMC_1692 D[1] Q[1] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_2 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_273 TSMC_274 TSMC_275 
+ TSMC_276 TSMC_1691 BWEB[2] TSMC_1692 D[2] Q[2] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_3 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_281 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_1691 BWEB[3] TSMC_1692 D[3] Q[3] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_4 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_289 TSMC_290 TSMC_291 
+ TSMC_292 TSMC_1691 BWEB[4] TSMC_1692 D[4] Q[4] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_5 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_297 TSMC_298 TSMC_299 
+ TSMC_300 TSMC_1691 BWEB[5] TSMC_1692 D[5] Q[5] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_6 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_305 TSMC_306 TSMC_307 
+ TSMC_308 TSMC_1691 BWEB[6] TSMC_1692 D[6] Q[6] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_7 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_313 TSMC_314 TSMC_315 
+ TSMC_316 TSMC_1691 BWEB[7] TSMC_1692 D[7] Q[7] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_8 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_321 TSMC_322 TSMC_323 
+ TSMC_324 TSMC_1691 BWEB[8] TSMC_1692 D[8] Q[8] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_9 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_329 TSMC_330 TSMC_331 
+ TSMC_332 TSMC_1691 BWEB[9] TSMC_1692 D[9] Q[9] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_10 TSMC_341 TSMC_342 TSMC_343 TSMC_344 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_1691 BWEB[10] TSMC_1692 D[10] Q[10] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_11 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_345 TSMC_346 TSMC_347 
+ TSMC_348 TSMC_1691 BWEB[11] TSMC_1692 D[11] Q[11] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_12 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_353 TSMC_354 TSMC_355 
+ TSMC_356 TSMC_1691 BWEB[12] TSMC_1692 D[12] Q[12] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_13 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_361 TSMC_362 TSMC_363 
+ TSMC_364 TSMC_1691 BWEB[13] TSMC_1692 D[13] Q[13] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_14 TSMC_373 TSMC_374 TSMC_375 TSMC_376 TSMC_369 TSMC_370 TSMC_371 
+ TSMC_372 TSMC_1691 BWEB[14] TSMC_1692 D[14] Q[14] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_L_15 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_377 TSMC_378 TSMC_379 
+ TSMC_380 TSMC_1691 BWEB[15] TSMC_1692 D[15] Q[15] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_16 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_385 TSMC_386 TSMC_387 
+ TSMC_388 TSMC_1702 BWEB[16] TSMC_1703 D[16] Q[16] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_17 TSMC_653 TSMC_654 TSMC_655 TSMC_656 TSMC_649 TSMC_650 TSMC_651 
+ TSMC_652 TSMC_1702 BWEB[17] TSMC_1703 D[17] Q[17] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_18 TSMC_661 TSMC_662 TSMC_663 TSMC_664 TSMC_657 TSMC_658 TSMC_659 
+ TSMC_660 TSMC_1702 BWEB[18] TSMC_1703 D[18] Q[18] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_19 TSMC_669 TSMC_670 TSMC_671 TSMC_672 TSMC_665 TSMC_666 TSMC_667 
+ TSMC_668 TSMC_1702 BWEB[19] TSMC_1703 D[19] Q[19] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_20 TSMC_677 TSMC_678 TSMC_679 TSMC_680 TSMC_673 TSMC_674 TSMC_675 
+ TSMC_676 TSMC_1702 BWEB[20] TSMC_1703 D[20] Q[20] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_21 TSMC_685 TSMC_686 TSMC_687 TSMC_688 TSMC_681 TSMC_682 TSMC_683 
+ TSMC_684 TSMC_1702 BWEB[21] TSMC_1703 D[21] Q[21] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_22 TSMC_693 TSMC_694 TSMC_695 TSMC_696 TSMC_689 TSMC_690 TSMC_691 
+ TSMC_692 TSMC_1702 BWEB[22] TSMC_1703 D[22] Q[22] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_23 TSMC_701 TSMC_702 TSMC_703 TSMC_704 TSMC_697 TSMC_698 TSMC_699 
+ TSMC_700 TSMC_1702 BWEB[23] TSMC_1703 D[23] Q[23] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_24 TSMC_709 TSMC_710 TSMC_711 TSMC_712 TSMC_705 TSMC_706 TSMC_707 
+ TSMC_708 TSMC_1702 BWEB[24] TSMC_1703 D[24] Q[24] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_25 TSMC_717 TSMC_718 TSMC_719 TSMC_720 TSMC_713 TSMC_714 TSMC_715 
+ TSMC_716 TSMC_1702 BWEB[25] TSMC_1703 D[25] Q[25] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_26 TSMC_725 TSMC_726 TSMC_727 TSMC_728 TSMC_721 TSMC_722 TSMC_723 
+ TSMC_724 TSMC_1702 BWEB[26] TSMC_1703 D[26] Q[26] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_27 TSMC_733 TSMC_734 TSMC_735 TSMC_736 TSMC_729 TSMC_730 TSMC_731 
+ TSMC_732 TSMC_1702 BWEB[27] TSMC_1703 D[27] Q[27] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_28 TSMC_741 TSMC_742 TSMC_743 TSMC_744 TSMC_737 TSMC_738 TSMC_739 
+ TSMC_740 TSMC_1702 BWEB[28] TSMC_1703 D[28] Q[28] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_29 TSMC_749 TSMC_750 TSMC_751 TSMC_752 TSMC_745 TSMC_746 TSMC_747 
+ TSMC_748 TSMC_1702 BWEB[29] TSMC_1703 D[29] Q[29] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_30 TSMC_757 TSMC_758 TSMC_759 TSMC_760 TSMC_753 TSMC_754 TSMC_755 
+ TSMC_756 TSMC_1702 BWEB[30] TSMC_1703 D[30] Q[30] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIOM4_R_31 TSMC_765 TSMC_766 TSMC_767 TSMC_768 TSMC_761 TSMC_762 TSMC_763 
+ TSMC_764 TSMC_1702 BWEB[31] TSMC_1703 D[31] Q[31] TSMC_1693 VDD VSS 
+ TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 
+ TSMC_1700 TSMC_1701 S1ALLSVTSW400W20_MIO_SB 
XMIO_SB_EDGE_L VDD TSMC_1704 TSMC_1705 VSS 
+ S1ALLSVTSW400W20_MIO_SB_EDGE 
XMIO_SB_EDGE_R VDD TSMC_1704 TSMC_1705 VSS 
+ S1ALLSVTSW400W20_MIO_SB_EDGE 
XCNT_M4_SB TSMC_1691 TSMC_1702 TSMC_1690 CEB TSMC_1692 TSMC_1703 CLK TSMC_771 
+ TSMC_772 TSMC_773 TSMC_774 TSMC_790 TSMC_791 TSMC_792 TSMC_793 
+ TSMC_779 TSMC_812 TSMC_841 TSMC_870 TSMC_899 TSMC_928 TSMC_957 
+ TSMC_986 TSMC_769 TSMC_1011 TSMC_1237 TSMC_1463 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 
+ TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 RTSEL[0] RTSEL[1] TSMC_1693 
+ TSMC_1705 TSMC_1689 VDD VSS WEB WTSEL[0] WTSEL[1] TSMC_1705 A[2] 
+ A[3] A[4] A[5] A[6] A[7] A[8] A[9] A[0] A[1] TSMC_1705 TSMC_1705 
+ S1ALLSVTSW400W20_CNT_M4_SB 
XD_WEB WEB TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_CEB CEB TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_CLK CLK TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A0 A[0] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A1 A[1] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A2 A[2] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A3 A[3] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A4 A[4] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A5 A[5] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A6 A[6] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A7 A[7] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A8 A[8] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_A9 A[9] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_D0 D[0] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D1 D[1] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D2 D[2] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D3 D[3] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D4 D[4] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D5 D[5] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D6 D[6] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D7 D[7] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D8 D[8] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D9 D[9] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D10 D[10] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D11 D[11] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D12 D[12] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D13 D[13] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D14 D[14] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D15 D[15] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D16 D[16] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D17 D[17] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D18 D[18] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D19 D[19] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D20 D[20] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D21 D[21] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D22 D[22] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D23 D[23] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D24 D[24] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D25 D[25] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D26 D[26] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D27 D[27] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D28 D[28] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D29 D[29] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D30 D[30] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_D31 D[31] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB0 BWEB[0] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB1 BWEB[1] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB2 BWEB[2] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB3 BWEB[3] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB4 BWEB[4] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB5 BWEB[5] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB6 BWEB[6] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB7 BWEB[7] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB8 BWEB[8] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB9 BWEB[9] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB10 BWEB[10] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB11 BWEB[11] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB12 BWEB[12] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB13 BWEB[13] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB14 BWEB[14] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB15 BWEB[15] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB16 BWEB[16] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB17 BWEB[17] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB18 BWEB[18] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB19 BWEB[19] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB20 BWEB[20] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB21 BWEB[21] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB22 BWEB[22] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB23 BWEB[23] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB24 BWEB[24] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB25 BWEB[25] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB26 BWEB[26] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB27 BWEB[27] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB28 BWEB[28] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB29 BWEB[29] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB30 BWEB[30] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_BWEB31 BWEB[31] VSS S1ALLSVTSW400W20_DIO_TALL 
XD_WTESL_1 WTSEL[1] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_WTESL_0 WTSEL[0] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_RTESL_1 RTSEL[1] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
XD_RTESL_0 RTSEL[0] TSMC_1705 VSS S1ALLSVTSW400W20_DIODE 
.ENDS


