# Created by MC2 : Version 2013.12.00.f on 2025/06/18, 12:00:46

 
###############################################################################
#                                                    
#        Technology     : TSMC 16nm CMOS Logic FinFet (FFC) HKMG
#        Memory Type    : TSMC 16nm FFC Two Port Register File with d130 bit cell
#        Library Name   : ts6n16ffcllsvta64x32m4fw (user specify : ts6n16ffcllsvta64x32m4fw)
#        Library Version: 170a
#        Generated Time : 2025/06/18, 11:59:49
###############################################################################
# STATEMENT OF USE                                                             
#                                                                              
#  This information contains confidential and proprietary information of TSMC. 
# No part of this information may be reproduced, transmitted, transcribed,     
# stored in a retrieval system, or translated into any human or computer       
# language, in any form or by any means, electronic, mechanical, magnetic,     
# optical, chemical, manual, or otherwise, without the prior written permission
# of TSMC. This information was prepared for informational purpose and is for  
# use by TSMC's customers only. TSMC reserves the right to make changes in the 
# inforrmation at any time and without notice.                                 
###############################################################################
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
#                                                                              

MACRO TS6N16FFCLLSVTA64X32M4FW
	CLASS BLOCK ;
	FOREIGN TS6N16FFCLLSVTA64X32M4FW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 16.957 BY 112.800 ;
	SYMMETRY X Y ;
	PIN AA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 52.142 16.957 52.222 ;
			LAYER M2 ;
			RECT 16.709 52.142 16.957 52.222 ;
			LAYER M3 ;
			RECT 16.709 52.142 16.957 52.222 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[0]

	PIN AA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 52.370 16.957 52.450 ;
			LAYER M2 ;
			RECT 16.709 52.370 16.957 52.450 ;
			LAYER M3 ;
			RECT 16.709 52.370 16.957 52.450 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[1]

	PIN AA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 55.334 16.957 55.414 ;
			LAYER M2 ;
			RECT 16.709 55.334 16.957 55.414 ;
			LAYER M3 ;
			RECT 16.709 55.334 16.957 55.414 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[2]

	PIN AA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 53.738 16.957 53.818 ;
			LAYER M2 ;
			RECT 16.709 53.738 16.957 53.818 ;
			LAYER M3 ;
			RECT 16.709 53.738 16.957 53.818 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[3]

	PIN AA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 55.106 16.957 55.186 ;
			LAYER M2 ;
			RECT 16.709 55.106 16.957 55.186 ;
			LAYER M3 ;
			RECT 16.709 55.106 16.957 55.186 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[4]

	PIN AA[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 53.966 16.957 54.046 ;
			LAYER M2 ;
			RECT 16.709 53.966 16.957 54.046 ;
			LAYER M3 ;
			RECT 16.709 53.966 16.957 54.046 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[5]

	PIN AB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 60.578 16.957 60.658 ;
			LAYER M2 ;
			RECT 16.709 60.578 16.957 60.658 ;
			LAYER M3 ;
			RECT 16.709 60.578 16.957 60.658 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[0]

	PIN AB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 60.350 16.957 60.430 ;
			LAYER M2 ;
			RECT 16.709 60.350 16.957 60.430 ;
			LAYER M3 ;
			RECT 16.709 60.350 16.957 60.430 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[1]

	PIN AB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 57.386 16.957 57.466 ;
			LAYER M2 ;
			RECT 16.709 57.386 16.957 57.466 ;
			LAYER M3 ;
			RECT 16.709 57.386 16.957 57.466 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[2]

	PIN AB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 58.982 16.957 59.062 ;
			LAYER M2 ;
			RECT 16.709 58.982 16.957 59.062 ;
			LAYER M3 ;
			RECT 16.709 58.982 16.957 59.062 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[3]

	PIN AB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 57.614 16.957 57.694 ;
			LAYER M2 ;
			RECT 16.709 57.614 16.957 57.694 ;
			LAYER M3 ;
			RECT 16.709 57.614 16.957 57.694 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[4]

	PIN AB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 58.754 16.957 58.834 ;
			LAYER M2 ;
			RECT 16.709 58.754 16.957 58.834 ;
			LAYER M3 ;
			RECT 16.709 58.754 16.957 58.834 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[5]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 1.799 16.957 1.879 ;
			LAYER M2 ;
			RECT 16.709 1.799 16.957 1.879 ;
			LAYER M3 ;
			RECT 16.709 1.799 16.957 1.879 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 4.679 16.957 4.759 ;
			LAYER M2 ;
			RECT 16.709 4.679 16.957 4.759 ;
			LAYER M3 ;
			RECT 16.709 4.679 16.957 4.759 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 7.559 16.957 7.639 ;
			LAYER M2 ;
			RECT 16.709 7.559 16.957 7.639 ;
			LAYER M3 ;
			RECT 16.709 7.559 16.957 7.639 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 10.439 16.957 10.519 ;
			LAYER M2 ;
			RECT 16.709 10.439 16.957 10.519 ;
			LAYER M3 ;
			RECT 16.709 10.439 16.957 10.519 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 13.319 16.957 13.399 ;
			LAYER M2 ;
			RECT 16.709 13.319 16.957 13.399 ;
			LAYER M3 ;
			RECT 16.709 13.319 16.957 13.399 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 16.199 16.957 16.279 ;
			LAYER M2 ;
			RECT 16.709 16.199 16.957 16.279 ;
			LAYER M3 ;
			RECT 16.709 16.199 16.957 16.279 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 19.079 16.957 19.159 ;
			LAYER M2 ;
			RECT 16.709 19.079 16.957 19.159 ;
			LAYER M3 ;
			RECT 16.709 19.079 16.957 19.159 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 21.959 16.957 22.039 ;
			LAYER M2 ;
			RECT 16.709 21.959 16.957 22.039 ;
			LAYER M3 ;
			RECT 16.709 21.959 16.957 22.039 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 24.839 16.957 24.919 ;
			LAYER M2 ;
			RECT 16.709 24.839 16.957 24.919 ;
			LAYER M3 ;
			RECT 16.709 24.839 16.957 24.919 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 27.719 16.957 27.799 ;
			LAYER M2 ;
			RECT 16.709 27.719 16.957 27.799 ;
			LAYER M3 ;
			RECT 16.709 27.719 16.957 27.799 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 30.599 16.957 30.679 ;
			LAYER M2 ;
			RECT 16.709 30.599 16.957 30.679 ;
			LAYER M3 ;
			RECT 16.709 30.599 16.957 30.679 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 33.479 16.957 33.559 ;
			LAYER M2 ;
			RECT 16.709 33.479 16.957 33.559 ;
			LAYER M3 ;
			RECT 16.709 33.479 16.957 33.559 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 36.359 16.957 36.439 ;
			LAYER M2 ;
			RECT 16.709 36.359 16.957 36.439 ;
			LAYER M3 ;
			RECT 16.709 36.359 16.957 36.439 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 39.239 16.957 39.319 ;
			LAYER M2 ;
			RECT 16.709 39.239 16.957 39.319 ;
			LAYER M3 ;
			RECT 16.709 39.239 16.957 39.319 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 42.119 16.957 42.199 ;
			LAYER M2 ;
			RECT 16.709 42.119 16.957 42.199 ;
			LAYER M3 ;
			RECT 16.709 42.119 16.957 42.199 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 44.999 16.957 45.079 ;
			LAYER M2 ;
			RECT 16.709 44.999 16.957 45.079 ;
			LAYER M3 ;
			RECT 16.709 44.999 16.957 45.079 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 67.721 16.957 67.801 ;
			LAYER M2 ;
			RECT 16.709 67.721 16.957 67.801 ;
			LAYER M3 ;
			RECT 16.709 67.721 16.957 67.801 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 70.601 16.957 70.681 ;
			LAYER M2 ;
			RECT 16.709 70.601 16.957 70.681 ;
			LAYER M3 ;
			RECT 16.709 70.601 16.957 70.681 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 73.481 16.957 73.561 ;
			LAYER M2 ;
			RECT 16.709 73.481 16.957 73.561 ;
			LAYER M3 ;
			RECT 16.709 73.481 16.957 73.561 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 76.361 16.957 76.441 ;
			LAYER M2 ;
			RECT 16.709 76.361 16.957 76.441 ;
			LAYER M3 ;
			RECT 16.709 76.361 16.957 76.441 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 79.241 16.957 79.321 ;
			LAYER M2 ;
			RECT 16.709 79.241 16.957 79.321 ;
			LAYER M3 ;
			RECT 16.709 79.241 16.957 79.321 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 82.121 16.957 82.201 ;
			LAYER M2 ;
			RECT 16.709 82.121 16.957 82.201 ;
			LAYER M3 ;
			RECT 16.709 82.121 16.957 82.201 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 85.001 16.957 85.081 ;
			LAYER M2 ;
			RECT 16.709 85.001 16.957 85.081 ;
			LAYER M3 ;
			RECT 16.709 85.001 16.957 85.081 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 87.881 16.957 87.961 ;
			LAYER M2 ;
			RECT 16.709 87.881 16.957 87.961 ;
			LAYER M3 ;
			RECT 16.709 87.881 16.957 87.961 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 90.761 16.957 90.841 ;
			LAYER M2 ;
			RECT 16.709 90.761 16.957 90.841 ;
			LAYER M3 ;
			RECT 16.709 90.761 16.957 90.841 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 93.641 16.957 93.721 ;
			LAYER M2 ;
			RECT 16.709 93.641 16.957 93.721 ;
			LAYER M3 ;
			RECT 16.709 93.641 16.957 93.721 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 96.521 16.957 96.601 ;
			LAYER M2 ;
			RECT 16.709 96.521 16.957 96.601 ;
			LAYER M3 ;
			RECT 16.709 96.521 16.957 96.601 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 99.401 16.957 99.481 ;
			LAYER M2 ;
			RECT 16.709 99.401 16.957 99.481 ;
			LAYER M3 ;
			RECT 16.709 99.401 16.957 99.481 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 102.281 16.957 102.361 ;
			LAYER M2 ;
			RECT 16.709 102.281 16.957 102.361 ;
			LAYER M3 ;
			RECT 16.709 102.281 16.957 102.361 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 105.161 16.957 105.241 ;
			LAYER M2 ;
			RECT 16.709 105.161 16.957 105.241 ;
			LAYER M3 ;
			RECT 16.709 105.161 16.957 105.241 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 108.041 16.957 108.121 ;
			LAYER M2 ;
			RECT 16.709 108.041 16.957 108.121 ;
			LAYER M3 ;
			RECT 16.709 108.041 16.957 108.121 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 110.921 16.957 111.001 ;
			LAYER M2 ;
			RECT 16.709 110.921 16.957 111.001 ;
			LAYER M3 ;
			RECT 16.709 110.921 16.957 111.001 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[31]

	PIN CLKR
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 63.314 16.957 63.394 ;
			LAYER M2 ;
			RECT 16.709 63.314 16.957 63.394 ;
			LAYER M3 ;
			RECT 16.709 63.314 16.957 63.394 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2280 LAYER M2 ;
		ANTENNAMAXAREACAR 40.1766 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0128 LAYER M3 ;
		ANTENNAMAXAREACAR 179.9160 LAYER M3 ;
	END CLKR

	PIN CLKW
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 48.722 16.957 48.802 ;
			LAYER M2 ;
			RECT 16.709 48.722 16.957 48.802 ;
			LAYER M3 ;
			RECT 16.709 48.722 16.957 48.802 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.4639 LAYER M2 ;
		ANTENNAMAXAREACAR 44.8112 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0082 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0159 LAYER M3 ;
		ANTENNAMAXAREACAR 150.9920 LAYER M3 ;
	END CLKW

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 2.951 16.957 3.031 ;
			LAYER M2 ;
			RECT 16.709 2.951 16.957 3.031 ;
			LAYER M3 ;
			RECT 16.709 2.951 16.957 3.031 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 5.831 16.957 5.911 ;
			LAYER M2 ;
			RECT 16.709 5.831 16.957 5.911 ;
			LAYER M3 ;
			RECT 16.709 5.831 16.957 5.911 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 8.711 16.957 8.791 ;
			LAYER M2 ;
			RECT 16.709 8.711 16.957 8.791 ;
			LAYER M3 ;
			RECT 16.709 8.711 16.957 8.791 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 11.591 16.957 11.671 ;
			LAYER M2 ;
			RECT 16.709 11.591 16.957 11.671 ;
			LAYER M3 ;
			RECT 16.709 11.591 16.957 11.671 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 14.471 16.957 14.551 ;
			LAYER M2 ;
			RECT 16.709 14.471 16.957 14.551 ;
			LAYER M3 ;
			RECT 16.709 14.471 16.957 14.551 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 17.351 16.957 17.431 ;
			LAYER M2 ;
			RECT 16.709 17.351 16.957 17.431 ;
			LAYER M3 ;
			RECT 16.709 17.351 16.957 17.431 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 20.231 16.957 20.311 ;
			LAYER M2 ;
			RECT 16.709 20.231 16.957 20.311 ;
			LAYER M3 ;
			RECT 16.709 20.231 16.957 20.311 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 23.111 16.957 23.191 ;
			LAYER M2 ;
			RECT 16.709 23.111 16.957 23.191 ;
			LAYER M3 ;
			RECT 16.709 23.111 16.957 23.191 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 25.991 16.957 26.071 ;
			LAYER M2 ;
			RECT 16.709 25.991 16.957 26.071 ;
			LAYER M3 ;
			RECT 16.709 25.991 16.957 26.071 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 28.871 16.957 28.951 ;
			LAYER M2 ;
			RECT 16.709 28.871 16.957 28.951 ;
			LAYER M3 ;
			RECT 16.709 28.871 16.957 28.951 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 31.751 16.957 31.831 ;
			LAYER M2 ;
			RECT 16.709 31.751 16.957 31.831 ;
			LAYER M3 ;
			RECT 16.709 31.751 16.957 31.831 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 34.631 16.957 34.711 ;
			LAYER M2 ;
			RECT 16.709 34.631 16.957 34.711 ;
			LAYER M3 ;
			RECT 16.709 34.631 16.957 34.711 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 37.511 16.957 37.591 ;
			LAYER M2 ;
			RECT 16.709 37.511 16.957 37.591 ;
			LAYER M3 ;
			RECT 16.709 37.511 16.957 37.591 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 40.391 16.957 40.471 ;
			LAYER M2 ;
			RECT 16.709 40.391 16.957 40.471 ;
			LAYER M3 ;
			RECT 16.709 40.391 16.957 40.471 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 43.271 16.957 43.351 ;
			LAYER M2 ;
			RECT 16.709 43.271 16.957 43.351 ;
			LAYER M3 ;
			RECT 16.709 43.271 16.957 43.351 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 46.151 16.957 46.231 ;
			LAYER M2 ;
			RECT 16.709 46.151 16.957 46.231 ;
			LAYER M3 ;
			RECT 16.709 46.151 16.957 46.231 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 66.569 16.957 66.649 ;
			LAYER M2 ;
			RECT 16.709 66.569 16.957 66.649 ;
			LAYER M3 ;
			RECT 16.709 66.569 16.957 66.649 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 69.449 16.957 69.529 ;
			LAYER M2 ;
			RECT 16.709 69.449 16.957 69.529 ;
			LAYER M3 ;
			RECT 16.709 69.449 16.957 69.529 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 72.329 16.957 72.409 ;
			LAYER M2 ;
			RECT 16.709 72.329 16.957 72.409 ;
			LAYER M3 ;
			RECT 16.709 72.329 16.957 72.409 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 75.209 16.957 75.289 ;
			LAYER M2 ;
			RECT 16.709 75.209 16.957 75.289 ;
			LAYER M3 ;
			RECT 16.709 75.209 16.957 75.289 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 78.089 16.957 78.169 ;
			LAYER M2 ;
			RECT 16.709 78.089 16.957 78.169 ;
			LAYER M3 ;
			RECT 16.709 78.089 16.957 78.169 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 80.969 16.957 81.049 ;
			LAYER M2 ;
			RECT 16.709 80.969 16.957 81.049 ;
			LAYER M3 ;
			RECT 16.709 80.969 16.957 81.049 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 83.849 16.957 83.929 ;
			LAYER M2 ;
			RECT 16.709 83.849 16.957 83.929 ;
			LAYER M3 ;
			RECT 16.709 83.849 16.957 83.929 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 86.729 16.957 86.809 ;
			LAYER M2 ;
			RECT 16.709 86.729 16.957 86.809 ;
			LAYER M3 ;
			RECT 16.709 86.729 16.957 86.809 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 89.609 16.957 89.689 ;
			LAYER M2 ;
			RECT 16.709 89.609 16.957 89.689 ;
			LAYER M3 ;
			RECT 16.709 89.609 16.957 89.689 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 92.489 16.957 92.569 ;
			LAYER M2 ;
			RECT 16.709 92.489 16.957 92.569 ;
			LAYER M3 ;
			RECT 16.709 92.489 16.957 92.569 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 95.369 16.957 95.449 ;
			LAYER M2 ;
			RECT 16.709 95.369 16.957 95.449 ;
			LAYER M3 ;
			RECT 16.709 95.369 16.957 95.449 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 98.249 16.957 98.329 ;
			LAYER M2 ;
			RECT 16.709 98.249 16.957 98.329 ;
			LAYER M3 ;
			RECT 16.709 98.249 16.957 98.329 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 101.129 16.957 101.209 ;
			LAYER M2 ;
			RECT 16.709 101.129 16.957 101.209 ;
			LAYER M3 ;
			RECT 16.709 101.129 16.957 101.209 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 104.009 16.957 104.089 ;
			LAYER M2 ;
			RECT 16.709 104.009 16.957 104.089 ;
			LAYER M3 ;
			RECT 16.709 104.009 16.957 104.089 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 106.889 16.957 106.969 ;
			LAYER M2 ;
			RECT 16.709 106.889 16.957 106.969 ;
			LAYER M3 ;
			RECT 16.709 106.889 16.957 106.969 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 109.769 16.957 109.849 ;
			LAYER M2 ;
			RECT 16.709 109.769 16.957 109.849 ;
			LAYER M3 ;
			RECT 16.709 109.769 16.957 109.849 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[31]

	PIN KP[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 50.090 16.957 50.170 ;
			LAYER M2 ;
			RECT 16.709 50.090 16.957 50.170 ;
			LAYER M3 ;
			RECT 16.709 50.090 16.957 50.170 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[0]

	PIN KP[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 50.318 16.957 50.398 ;
			LAYER M2 ;
			RECT 16.709 50.318 16.957 50.398 ;
			LAYER M3 ;
			RECT 16.709 50.318 16.957 50.398 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[1]

	PIN KP[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 50.546 16.957 50.626 ;
			LAYER M2 ;
			RECT 16.709 50.546 16.957 50.626 ;
			LAYER M3 ;
			RECT 16.709 50.546 16.957 50.626 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[2]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 2.375 16.957 2.455 ;
			LAYER M2 ;
			RECT 16.709 2.375 16.957 2.455 ;
			LAYER M3 ;
			RECT 16.709 2.375 16.957 2.455 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 5.255 16.957 5.335 ;
			LAYER M2 ;
			RECT 16.709 5.255 16.957 5.335 ;
			LAYER M3 ;
			RECT 16.709 5.255 16.957 5.335 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 8.135 16.957 8.215 ;
			LAYER M2 ;
			RECT 16.709 8.135 16.957 8.215 ;
			LAYER M3 ;
			RECT 16.709 8.135 16.957 8.215 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 11.015 16.957 11.095 ;
			LAYER M2 ;
			RECT 16.709 11.015 16.957 11.095 ;
			LAYER M3 ;
			RECT 16.709 11.015 16.957 11.095 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 13.895 16.957 13.975 ;
			LAYER M2 ;
			RECT 16.709 13.895 16.957 13.975 ;
			LAYER M3 ;
			RECT 16.709 13.895 16.957 13.975 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 16.775 16.957 16.855 ;
			LAYER M2 ;
			RECT 16.709 16.775 16.957 16.855 ;
			LAYER M3 ;
			RECT 16.709 16.775 16.957 16.855 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 19.655 16.957 19.735 ;
			LAYER M2 ;
			RECT 16.709 19.655 16.957 19.735 ;
			LAYER M3 ;
			RECT 16.709 19.655 16.957 19.735 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 22.535 16.957 22.615 ;
			LAYER M2 ;
			RECT 16.709 22.535 16.957 22.615 ;
			LAYER M3 ;
			RECT 16.709 22.535 16.957 22.615 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 25.415 16.957 25.495 ;
			LAYER M2 ;
			RECT 16.709 25.415 16.957 25.495 ;
			LAYER M3 ;
			RECT 16.709 25.415 16.957 25.495 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 28.295 16.957 28.375 ;
			LAYER M2 ;
			RECT 16.709 28.295 16.957 28.375 ;
			LAYER M3 ;
			RECT 16.709 28.295 16.957 28.375 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 31.175 16.957 31.255 ;
			LAYER M2 ;
			RECT 16.709 31.175 16.957 31.255 ;
			LAYER M3 ;
			RECT 16.709 31.175 16.957 31.255 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 34.055 16.957 34.135 ;
			LAYER M2 ;
			RECT 16.709 34.055 16.957 34.135 ;
			LAYER M3 ;
			RECT 16.709 34.055 16.957 34.135 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 36.935 16.957 37.015 ;
			LAYER M2 ;
			RECT 16.709 36.935 16.957 37.015 ;
			LAYER M3 ;
			RECT 16.709 36.935 16.957 37.015 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 39.815 16.957 39.895 ;
			LAYER M2 ;
			RECT 16.709 39.815 16.957 39.895 ;
			LAYER M3 ;
			RECT 16.709 39.815 16.957 39.895 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 42.695 16.957 42.775 ;
			LAYER M2 ;
			RECT 16.709 42.695 16.957 42.775 ;
			LAYER M3 ;
			RECT 16.709 42.695 16.957 42.775 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 45.575 16.957 45.655 ;
			LAYER M2 ;
			RECT 16.709 45.575 16.957 45.655 ;
			LAYER M3 ;
			RECT 16.709 45.575 16.957 45.655 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 67.145 16.957 67.225 ;
			LAYER M2 ;
			RECT 16.709 67.145 16.957 67.225 ;
			LAYER M3 ;
			RECT 16.709 67.145 16.957 67.225 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 70.025 16.957 70.105 ;
			LAYER M2 ;
			RECT 16.709 70.025 16.957 70.105 ;
			LAYER M3 ;
			RECT 16.709 70.025 16.957 70.105 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 72.905 16.957 72.985 ;
			LAYER M2 ;
			RECT 16.709 72.905 16.957 72.985 ;
			LAYER M3 ;
			RECT 16.709 72.905 16.957 72.985 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 75.785 16.957 75.865 ;
			LAYER M2 ;
			RECT 16.709 75.785 16.957 75.865 ;
			LAYER M3 ;
			RECT 16.709 75.785 16.957 75.865 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 78.665 16.957 78.745 ;
			LAYER M2 ;
			RECT 16.709 78.665 16.957 78.745 ;
			LAYER M3 ;
			RECT 16.709 78.665 16.957 78.745 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 81.545 16.957 81.625 ;
			LAYER M2 ;
			RECT 16.709 81.545 16.957 81.625 ;
			LAYER M3 ;
			RECT 16.709 81.545 16.957 81.625 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 84.425 16.957 84.505 ;
			LAYER M2 ;
			RECT 16.709 84.425 16.957 84.505 ;
			LAYER M3 ;
			RECT 16.709 84.425 16.957 84.505 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 87.305 16.957 87.385 ;
			LAYER M2 ;
			RECT 16.709 87.305 16.957 87.385 ;
			LAYER M3 ;
			RECT 16.709 87.305 16.957 87.385 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 90.185 16.957 90.265 ;
			LAYER M2 ;
			RECT 16.709 90.185 16.957 90.265 ;
			LAYER M3 ;
			RECT 16.709 90.185 16.957 90.265 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 93.065 16.957 93.145 ;
			LAYER M2 ;
			RECT 16.709 93.065 16.957 93.145 ;
			LAYER M3 ;
			RECT 16.709 93.065 16.957 93.145 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 95.945 16.957 96.025 ;
			LAYER M2 ;
			RECT 16.709 95.945 16.957 96.025 ;
			LAYER M3 ;
			RECT 16.709 95.945 16.957 96.025 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 98.825 16.957 98.905 ;
			LAYER M2 ;
			RECT 16.709 98.825 16.957 98.905 ;
			LAYER M3 ;
			RECT 16.709 98.825 16.957 98.905 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 101.705 16.957 101.785 ;
			LAYER M2 ;
			RECT 16.709 101.705 16.957 101.785 ;
			LAYER M3 ;
			RECT 16.709 101.705 16.957 101.785 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 104.585 16.957 104.665 ;
			LAYER M2 ;
			RECT 16.709 104.585 16.957 104.665 ;
			LAYER M3 ;
			RECT 16.709 104.585 16.957 104.665 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 107.465 16.957 107.545 ;
			LAYER M2 ;
			RECT 16.709 107.465 16.957 107.545 ;
			LAYER M3 ;
			RECT 16.709 107.465 16.957 107.545 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 110.345 16.957 110.425 ;
			LAYER M2 ;
			RECT 16.709 110.345 16.957 110.425 ;
			LAYER M3 ;
			RECT 16.709 110.345 16.957 110.425 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[31]

	PIN RCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 65.138 16.957 65.218 ;
			LAYER M2 ;
			RECT 16.709 65.138 16.957 65.218 ;
			LAYER M3 ;
			RECT 16.709 65.138 16.957 65.218 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[0]

	PIN RCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 64.910 16.957 64.990 ;
			LAYER M2 ;
			RECT 16.709 64.910 16.957 64.990 ;
			LAYER M3 ;
			RECT 16.709 64.910 16.957 64.990 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[1]

	PIN REB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 61.490 16.957 61.570 ;
			LAYER M2 ;
			RECT 16.709 61.490 16.957 61.570 ;
			LAYER M3 ;
			RECT 16.709 61.490 16.957 61.570 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0860 LAYER M1 ;
		ANTENNAMAXAREACAR 12.8828 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0840 LAYER M2 ;
		ANTENNAMAXAREACAR 20.5069 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4602 LAYER M3 ;
		ANTENNAMAXAREACAR 218.8550 LAYER M3 ;
	END REB

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.624 16.837 1.784 ;
			LAYER M4 ;
			RECT 0.120 3.064 16.837 3.224 ;
			LAYER M4 ;
			RECT 0.120 4.504 16.837 4.664 ;
			LAYER M4 ;
			RECT 0.120 5.944 16.837 6.104 ;
			LAYER M4 ;
			RECT 0.120 7.384 16.837 7.544 ;
			LAYER M4 ;
			RECT 0.120 8.824 16.837 8.984 ;
			LAYER M4 ;
			RECT 0.120 10.264 16.837 10.424 ;
			LAYER M4 ;
			RECT 0.120 11.704 16.837 11.864 ;
			LAYER M4 ;
			RECT 0.120 13.144 16.837 13.304 ;
			LAYER M4 ;
			RECT 0.120 14.584 16.837 14.744 ;
			LAYER M4 ;
			RECT 0.120 16.024 16.837 16.184 ;
			LAYER M4 ;
			RECT 0.120 17.464 16.837 17.624 ;
			LAYER M4 ;
			RECT 0.120 18.904 16.837 19.064 ;
			LAYER M4 ;
			RECT 0.120 20.344 16.837 20.504 ;
			LAYER M4 ;
			RECT 0.120 21.784 16.837 21.944 ;
			LAYER M4 ;
			RECT 0.120 23.224 16.837 23.384 ;
			LAYER M4 ;
			RECT 0.120 24.664 16.837 24.824 ;
			LAYER M4 ;
			RECT 0.120 26.104 16.837 26.264 ;
			LAYER M4 ;
			RECT 0.120 27.544 16.837 27.704 ;
			LAYER M4 ;
			RECT 0.120 28.984 16.837 29.144 ;
			LAYER M4 ;
			RECT 0.120 30.424 16.837 30.584 ;
			LAYER M4 ;
			RECT 0.120 31.864 16.837 32.024 ;
			LAYER M4 ;
			RECT 0.120 33.304 16.837 33.464 ;
			LAYER M4 ;
			RECT 0.120 34.744 16.837 34.904 ;
			LAYER M4 ;
			RECT 0.120 36.184 16.837 36.344 ;
			LAYER M4 ;
			RECT 0.120 37.624 16.837 37.784 ;
			LAYER M4 ;
			RECT 0.120 39.064 16.837 39.224 ;
			LAYER M4 ;
			RECT 0.120 40.504 16.837 40.664 ;
			LAYER M4 ;
			RECT 0.120 41.944 16.837 42.104 ;
			LAYER M4 ;
			RECT 0.120 43.384 16.837 43.544 ;
			LAYER M4 ;
			RECT 0.120 44.824 16.837 44.984 ;
			LAYER M4 ;
			RECT 0.120 46.264 16.837 46.424 ;
			LAYER M4 ;
			RECT 0.120 47.684 16.837 47.884 ;
			LAYER M4 ;
			RECT 0.120 48.620 16.837 48.820 ;
			LAYER M4 ;
			RECT 0.120 50.156 16.837 50.356 ;
			LAYER M4 ;
			RECT 0.120 51.692 16.837 51.892 ;
			LAYER M4 ;
			RECT 0.120 53.228 16.837 53.428 ;
			LAYER M4 ;
			RECT 0.120 54.764 16.837 54.964 ;
			LAYER M4 ;
			RECT 0.120 56.300 16.837 56.500 ;
			LAYER M4 ;
			RECT 0.120 57.836 16.837 58.036 ;
			LAYER M4 ;
			RECT 0.120 59.372 16.837 59.572 ;
			LAYER M4 ;
			RECT 0.120 60.908 16.837 61.108 ;
			LAYER M4 ;
			RECT 0.120 62.444 16.837 62.644 ;
			LAYER M4 ;
			RECT 0.120 63.980 16.837 64.180 ;
			LAYER M4 ;
			RECT 0.120 64.916 16.837 65.116 ;
			LAYER M4 ;
			RECT 0.120 66.376 16.837 66.536 ;
			LAYER M4 ;
			RECT 0.120 67.816 16.837 67.976 ;
			LAYER M4 ;
			RECT 0.120 69.256 16.837 69.416 ;
			LAYER M4 ;
			RECT 0.120 70.696 16.837 70.856 ;
			LAYER M4 ;
			RECT 0.120 72.136 16.837 72.296 ;
			LAYER M4 ;
			RECT 0.120 73.576 16.837 73.736 ;
			LAYER M4 ;
			RECT 0.120 75.016 16.837 75.176 ;
			LAYER M4 ;
			RECT 0.120 76.456 16.837 76.616 ;
			LAYER M4 ;
			RECT 0.120 77.896 16.837 78.056 ;
			LAYER M4 ;
			RECT 0.120 79.336 16.837 79.496 ;
			LAYER M4 ;
			RECT 0.120 80.776 16.837 80.936 ;
			LAYER M4 ;
			RECT 0.120 82.216 16.837 82.376 ;
			LAYER M4 ;
			RECT 0.120 83.656 16.837 83.816 ;
			LAYER M4 ;
			RECT 0.120 85.096 16.837 85.256 ;
			LAYER M4 ;
			RECT 0.120 86.536 16.837 86.696 ;
			LAYER M4 ;
			RECT 0.120 87.976 16.837 88.136 ;
			LAYER M4 ;
			RECT 0.120 89.416 16.837 89.576 ;
			LAYER M4 ;
			RECT 0.120 90.856 16.837 91.016 ;
			LAYER M4 ;
			RECT 0.120 92.296 16.837 92.456 ;
			LAYER M4 ;
			RECT 0.120 93.736 16.837 93.896 ;
			LAYER M4 ;
			RECT 0.120 95.176 16.837 95.336 ;
			LAYER M4 ;
			RECT 0.120 96.616 16.837 96.776 ;
			LAYER M4 ;
			RECT 0.120 98.056 16.837 98.216 ;
			LAYER M4 ;
			RECT 0.120 99.496 16.837 99.656 ;
			LAYER M4 ;
			RECT 0.120 100.936 16.837 101.096 ;
			LAYER M4 ;
			RECT 0.120 102.376 16.837 102.536 ;
			LAYER M4 ;
			RECT 0.120 103.816 16.837 103.976 ;
			LAYER M4 ;
			RECT 0.120 105.256 16.837 105.416 ;
			LAYER M4 ;
			RECT 0.120 106.696 16.837 106.856 ;
			LAYER M4 ;
			RECT 0.120 108.136 16.837 108.296 ;
			LAYER M4 ;
			RECT 0.120 109.576 16.837 109.736 ;
			LAYER M4 ;
			RECT 0.120 111.016 16.837 111.176 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 0.884 16.837 1.084 ;
			LAYER M4 ;
			RECT 0.120 2.324 16.837 2.524 ;
			LAYER M4 ;
			RECT 0.120 3.764 16.837 3.964 ;
			LAYER M4 ;
			RECT 0.120 5.204 16.837 5.404 ;
			LAYER M4 ;
			RECT 0.120 6.644 16.837 6.844 ;
			LAYER M4 ;
			RECT 0.120 8.084 16.837 8.284 ;
			LAYER M4 ;
			RECT 0.120 9.524 16.837 9.724 ;
			LAYER M4 ;
			RECT 0.120 10.964 16.837 11.164 ;
			LAYER M4 ;
			RECT 0.120 12.404 16.837 12.604 ;
			LAYER M4 ;
			RECT 0.120 13.844 16.837 14.044 ;
			LAYER M4 ;
			RECT 0.120 15.284 16.837 15.484 ;
			LAYER M4 ;
			RECT 0.120 16.724 16.837 16.924 ;
			LAYER M4 ;
			RECT 0.120 18.164 16.837 18.364 ;
			LAYER M4 ;
			RECT 0.120 19.604 16.837 19.804 ;
			LAYER M4 ;
			RECT 0.120 21.044 16.837 21.244 ;
			LAYER M4 ;
			RECT 0.120 22.484 16.837 22.684 ;
			LAYER M4 ;
			RECT 0.120 23.924 16.837 24.124 ;
			LAYER M4 ;
			RECT 0.120 25.364 16.837 25.564 ;
			LAYER M4 ;
			RECT 0.120 26.804 16.837 27.004 ;
			LAYER M4 ;
			RECT 0.120 28.244 16.837 28.444 ;
			LAYER M4 ;
			RECT 0.120 29.684 16.837 29.884 ;
			LAYER M4 ;
			RECT 0.120 31.124 16.837 31.324 ;
			LAYER M4 ;
			RECT 0.120 32.564 16.837 32.764 ;
			LAYER M4 ;
			RECT 0.120 34.004 16.837 34.204 ;
			LAYER M4 ;
			RECT 0.120 35.444 16.837 35.644 ;
			LAYER M4 ;
			RECT 0.120 36.884 16.837 37.084 ;
			LAYER M4 ;
			RECT 0.120 38.324 16.837 38.524 ;
			LAYER M4 ;
			RECT 0.120 39.764 16.837 39.964 ;
			LAYER M4 ;
			RECT 0.120 41.204 16.837 41.404 ;
			LAYER M4 ;
			RECT 0.120 42.644 16.837 42.844 ;
			LAYER M4 ;
			RECT 0.120 44.084 16.837 44.284 ;
			LAYER M4 ;
			RECT 0.120 45.524 16.837 45.724 ;
			LAYER M4 ;
			RECT 0.120 46.964 16.837 47.164 ;
			LAYER M4 ;
			RECT 0.120 49.388 16.837 49.588 ;
			LAYER M4 ;
			RECT 0.120 50.924 16.837 51.124 ;
			LAYER M4 ;
			RECT 0.120 52.460 16.837 52.660 ;
			LAYER M4 ;
			RECT 0.120 53.996 16.837 54.196 ;
			LAYER M4 ;
			RECT 0.120 55.532 16.837 55.732 ;
			LAYER M4 ;
			RECT 0.120 57.068 16.837 57.268 ;
			LAYER M4 ;
			RECT 0.120 58.604 16.837 58.804 ;
			LAYER M4 ;
			RECT 0.120 60.140 16.837 60.340 ;
			LAYER M4 ;
			RECT 0.120 61.676 16.837 61.876 ;
			LAYER M4 ;
			RECT 0.120 63.212 16.837 63.412 ;
			LAYER M4 ;
			RECT 0.120 65.636 16.837 65.836 ;
			LAYER M4 ;
			RECT 0.120 67.076 16.837 67.276 ;
			LAYER M4 ;
			RECT 0.120 68.516 16.837 68.716 ;
			LAYER M4 ;
			RECT 0.120 69.956 16.837 70.156 ;
			LAYER M4 ;
			RECT 0.120 71.396 16.837 71.596 ;
			LAYER M4 ;
			RECT 0.120 72.836 16.837 73.036 ;
			LAYER M4 ;
			RECT 0.120 74.276 16.837 74.476 ;
			LAYER M4 ;
			RECT 0.120 75.716 16.837 75.916 ;
			LAYER M4 ;
			RECT 0.120 77.156 16.837 77.356 ;
			LAYER M4 ;
			RECT 0.120 78.596 16.837 78.796 ;
			LAYER M4 ;
			RECT 0.120 80.036 16.837 80.236 ;
			LAYER M4 ;
			RECT 0.120 81.476 16.837 81.676 ;
			LAYER M4 ;
			RECT 0.120 82.916 16.837 83.116 ;
			LAYER M4 ;
			RECT 0.120 84.356 16.837 84.556 ;
			LAYER M4 ;
			RECT 0.120 85.796 16.837 85.996 ;
			LAYER M4 ;
			RECT 0.120 87.236 16.837 87.436 ;
			LAYER M4 ;
			RECT 0.120 88.676 16.837 88.876 ;
			LAYER M4 ;
			RECT 0.120 90.116 16.837 90.316 ;
			LAYER M4 ;
			RECT 0.120 91.556 16.837 91.756 ;
			LAYER M4 ;
			RECT 0.120 92.996 16.837 93.196 ;
			LAYER M4 ;
			RECT 0.120 94.436 16.837 94.636 ;
			LAYER M4 ;
			RECT 0.120 95.876 16.837 96.076 ;
			LAYER M4 ;
			RECT 0.120 97.316 16.837 97.516 ;
			LAYER M4 ;
			RECT 0.120 98.756 16.837 98.956 ;
			LAYER M4 ;
			RECT 0.120 100.196 16.837 100.396 ;
			LAYER M4 ;
			RECT 0.120 101.636 16.837 101.836 ;
			LAYER M4 ;
			RECT 0.120 103.076 16.837 103.276 ;
			LAYER M4 ;
			RECT 0.120 104.516 16.837 104.716 ;
			LAYER M4 ;
			RECT 0.120 105.956 16.837 106.156 ;
			LAYER M4 ;
			RECT 0.120 107.396 16.837 107.596 ;
			LAYER M4 ;
			RECT 0.120 108.836 16.837 109.036 ;
			LAYER M4 ;
			RECT 0.120 110.276 16.837 110.476 ;
			LAYER M4 ;
			RECT 0.120 111.716 16.837 111.916 ;
		END
	END VSS

	PIN WCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 48.038 16.957 48.118 ;
			LAYER M2 ;
			RECT 16.709 48.038 16.957 48.118 ;
			LAYER M3 ;
			RECT 16.709 48.038 16.957 48.118 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[0]

	PIN WCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 47.810 16.957 47.890 ;
			LAYER M2 ;
			RECT 16.709 47.810 16.957 47.890 ;
			LAYER M3 ;
			RECT 16.709 47.810 16.957 47.890 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.709 51.230 16.957 51.310 ;
			LAYER M2 ;
			RECT 16.709 51.230 16.957 51.310 ;
			LAYER M3 ;
			RECT 16.709 51.230 16.957 51.310 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0886 LAYER M1 ;
		ANTENNAMAXAREACAR 9.6368 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0833 LAYER M2 ;
		ANTENNAMAXAREACAR 13.2425 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4593 LAYER M3 ;
		ANTENNAMAXAREACAR 211.0720 LAYER M3 ;
	END WEB

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 16.957 112.800 ;
		LAYER M2 ;
		RECT 0.000 0.000 16.957 112.800 ;
		LAYER M3 ;
		RECT 0.000 0.000 16.957 112.800 ;
		LAYER M4 ;
		RECT 0.227 0.524 16.407 0.724 ;
		LAYER M4 ;
		RECT 0.227 1.358 15.977 1.518 ;
		LAYER M4 ;
		RECT 0.227 1.890 15.977 2.050 ;
		LAYER M4 ;
		RECT 0.227 2.798 15.977 2.958 ;
		LAYER M4 ;
		RECT 0.227 3.330 15.977 3.490 ;
		LAYER M4 ;
		RECT 0.227 4.238 15.977 4.398 ;
		LAYER M4 ;
		RECT 0.227 4.770 15.977 4.930 ;
		LAYER M4 ;
		RECT 0.227 5.678 15.977 5.838 ;
		LAYER M4 ;
		RECT 0.227 6.210 15.977 6.370 ;
		LAYER M4 ;
		RECT 0.227 7.118 15.977 7.278 ;
		LAYER M4 ;
		RECT 0.227 7.650 15.977 7.810 ;
		LAYER M4 ;
		RECT 0.227 8.558 15.977 8.718 ;
		LAYER M4 ;
		RECT 0.227 9.090 15.977 9.250 ;
		LAYER M4 ;
		RECT 0.227 9.998 15.977 10.158 ;
		LAYER M4 ;
		RECT 0.227 10.530 15.977 10.690 ;
		LAYER M4 ;
		RECT 0.227 11.438 15.977 11.598 ;
		LAYER M4 ;
		RECT 0.227 11.970 15.977 12.130 ;
		LAYER M4 ;
		RECT 0.227 12.878 15.977 13.038 ;
		LAYER M4 ;
		RECT 0.227 13.410 15.977 13.570 ;
		LAYER M4 ;
		RECT 0.227 14.318 15.977 14.478 ;
		LAYER M4 ;
		RECT 0.227 14.850 15.977 15.010 ;
		LAYER M4 ;
		RECT 0.227 15.758 15.977 15.918 ;
		LAYER M4 ;
		RECT 0.227 16.290 15.977 16.450 ;
		LAYER M4 ;
		RECT 0.227 17.198 15.977 17.358 ;
		LAYER M4 ;
		RECT 0.227 17.730 15.977 17.890 ;
		LAYER M4 ;
		RECT 0.227 18.638 15.977 18.798 ;
		LAYER M4 ;
		RECT 0.227 19.170 15.977 19.330 ;
		LAYER M4 ;
		RECT 0.227 20.078 15.977 20.238 ;
		LAYER M4 ;
		RECT 0.227 20.610 15.977 20.770 ;
		LAYER M4 ;
		RECT 0.227 21.518 15.977 21.678 ;
		LAYER M4 ;
		RECT 0.227 22.050 15.977 22.210 ;
		LAYER M4 ;
		RECT 0.227 22.958 15.977 23.118 ;
		LAYER M4 ;
		RECT 0.227 23.490 15.977 23.650 ;
		LAYER M4 ;
		RECT 0.227 24.398 15.977 24.558 ;
		LAYER M4 ;
		RECT 0.227 24.930 15.977 25.090 ;
		LAYER M4 ;
		RECT 0.227 25.838 15.977 25.998 ;
		LAYER M4 ;
		RECT 0.227 26.370 15.977 26.530 ;
		LAYER M4 ;
		RECT 0.227 27.278 15.977 27.438 ;
		LAYER M4 ;
		RECT 0.227 27.810 15.977 27.970 ;
		LAYER M4 ;
		RECT 0.227 28.718 15.977 28.878 ;
		LAYER M4 ;
		RECT 0.227 29.250 15.977 29.410 ;
		LAYER M4 ;
		RECT 0.227 30.158 15.977 30.318 ;
		LAYER M4 ;
		RECT 0.227 30.690 15.977 30.850 ;
		LAYER M4 ;
		RECT 0.227 31.598 15.977 31.758 ;
		LAYER M4 ;
		RECT 0.227 32.130 15.977 32.290 ;
		LAYER M4 ;
		RECT 0.227 33.038 15.977 33.198 ;
		LAYER M4 ;
		RECT 0.227 33.570 15.977 33.730 ;
		LAYER M4 ;
		RECT 0.227 34.478 15.977 34.638 ;
		LAYER M4 ;
		RECT 0.227 35.010 15.977 35.170 ;
		LAYER M4 ;
		RECT 0.227 35.918 15.977 36.078 ;
		LAYER M4 ;
		RECT 0.227 36.450 15.977 36.610 ;
		LAYER M4 ;
		RECT 0.227 37.358 15.977 37.518 ;
		LAYER M4 ;
		RECT 0.227 37.890 15.977 38.050 ;
		LAYER M4 ;
		RECT 0.227 38.798 15.977 38.958 ;
		LAYER M4 ;
		RECT 0.227 39.330 15.977 39.490 ;
		LAYER M4 ;
		RECT 0.227 40.238 15.977 40.398 ;
		LAYER M4 ;
		RECT 0.227 40.770 15.977 40.930 ;
		LAYER M4 ;
		RECT 0.227 41.678 15.977 41.838 ;
		LAYER M4 ;
		RECT 0.227 42.210 15.977 42.370 ;
		LAYER M4 ;
		RECT 0.227 43.118 15.977 43.278 ;
		LAYER M4 ;
		RECT 0.227 43.650 15.977 43.810 ;
		LAYER M4 ;
		RECT 0.227 44.558 15.977 44.718 ;
		LAYER M4 ;
		RECT 0.227 45.090 15.977 45.250 ;
		LAYER M4 ;
		RECT 0.227 45.998 15.977 46.158 ;
		LAYER M4 ;
		RECT 0.227 46.530 15.977 46.690 ;
		LAYER M4 ;
		RECT 0.227 47.324 15.977 47.524 ;
		LAYER M4 ;
		RECT 0.227 48.236 15.977 48.436 ;
		LAYER M4 ;
		RECT 0.227 49.004 15.977 49.204 ;
		LAYER M4 ;
		RECT 0.227 49.772 15.977 49.972 ;
		LAYER M4 ;
		RECT 0.227 50.540 15.977 50.740 ;
		LAYER M4 ;
		RECT 0.227 51.308 15.977 51.508 ;
		LAYER M4 ;
		RECT 0.227 52.076 15.977 52.276 ;
		LAYER M4 ;
		RECT 0.227 52.844 15.977 53.044 ;
		LAYER M4 ;
		RECT 0.227 53.612 15.977 53.812 ;
		LAYER M4 ;
		RECT 0.227 54.380 15.977 54.580 ;
		LAYER M4 ;
		RECT 0.227 55.148 15.977 55.348 ;
		LAYER M4 ;
		RECT 0.227 55.916 15.977 56.116 ;
		LAYER M4 ;
		RECT 0.227 56.684 15.977 56.884 ;
		LAYER M4 ;
		RECT 0.227 57.452 15.977 57.652 ;
		LAYER M4 ;
		RECT 0.227 58.220 15.977 58.420 ;
		LAYER M4 ;
		RECT 0.227 58.988 15.977 59.188 ;
		LAYER M4 ;
		RECT 0.227 59.756 15.977 59.956 ;
		LAYER M4 ;
		RECT 0.227 60.524 15.977 60.724 ;
		LAYER M4 ;
		RECT 0.227 61.292 15.977 61.492 ;
		LAYER M4 ;
		RECT 0.227 62.060 15.977 62.260 ;
		LAYER M4 ;
		RECT 0.227 62.828 15.977 63.028 ;
		LAYER M4 ;
		RECT 0.227 63.596 15.977 63.796 ;
		LAYER M4 ;
		RECT 0.227 64.364 15.977 64.564 ;
		LAYER M4 ;
		RECT 0.227 65.276 15.977 65.476 ;
		LAYER M4 ;
		RECT 0.227 66.110 15.977 66.270 ;
		LAYER M4 ;
		RECT 0.227 66.642 15.977 66.802 ;
		LAYER M4 ;
		RECT 0.227 67.550 15.977 67.710 ;
		LAYER M4 ;
		RECT 0.227 68.082 15.977 68.242 ;
		LAYER M4 ;
		RECT 0.227 68.990 15.977 69.150 ;
		LAYER M4 ;
		RECT 0.227 69.522 15.977 69.682 ;
		LAYER M4 ;
		RECT 0.227 70.430 15.977 70.590 ;
		LAYER M4 ;
		RECT 0.227 70.962 15.977 71.122 ;
		LAYER M4 ;
		RECT 0.227 71.870 15.977 72.030 ;
		LAYER M4 ;
		RECT 0.227 72.402 15.977 72.562 ;
		LAYER M4 ;
		RECT 0.227 73.310 15.977 73.470 ;
		LAYER M4 ;
		RECT 0.227 73.842 15.977 74.002 ;
		LAYER M4 ;
		RECT 0.227 74.750 15.977 74.910 ;
		LAYER M4 ;
		RECT 0.227 75.282 15.977 75.442 ;
		LAYER M4 ;
		RECT 0.227 76.190 15.977 76.350 ;
		LAYER M4 ;
		RECT 0.227 76.722 15.977 76.882 ;
		LAYER M4 ;
		RECT 0.227 77.630 15.977 77.790 ;
		LAYER M4 ;
		RECT 0.227 78.162 15.977 78.322 ;
		LAYER M4 ;
		RECT 0.227 79.070 15.977 79.230 ;
		LAYER M4 ;
		RECT 0.227 79.602 15.977 79.762 ;
		LAYER M4 ;
		RECT 0.227 80.510 15.977 80.670 ;
		LAYER M4 ;
		RECT 0.227 81.042 15.977 81.202 ;
		LAYER M4 ;
		RECT 0.227 81.950 15.977 82.110 ;
		LAYER M4 ;
		RECT 0.227 82.482 15.977 82.642 ;
		LAYER M4 ;
		RECT 0.227 83.390 15.977 83.550 ;
		LAYER M4 ;
		RECT 0.227 83.922 15.977 84.082 ;
		LAYER M4 ;
		RECT 0.227 84.830 15.977 84.990 ;
		LAYER M4 ;
		RECT 0.227 85.362 15.977 85.522 ;
		LAYER M4 ;
		RECT 0.227 86.270 15.977 86.430 ;
		LAYER M4 ;
		RECT 0.227 86.802 15.977 86.962 ;
		LAYER M4 ;
		RECT 0.227 87.710 15.977 87.870 ;
		LAYER M4 ;
		RECT 0.227 88.242 15.977 88.402 ;
		LAYER M4 ;
		RECT 0.227 89.150 15.977 89.310 ;
		LAYER M4 ;
		RECT 0.227 89.682 15.977 89.842 ;
		LAYER M4 ;
		RECT 0.227 90.590 15.977 90.750 ;
		LAYER M4 ;
		RECT 0.227 91.122 15.977 91.282 ;
		LAYER M4 ;
		RECT 0.227 92.030 15.977 92.190 ;
		LAYER M4 ;
		RECT 0.227 92.562 15.977 92.722 ;
		LAYER M4 ;
		RECT 0.227 93.470 15.977 93.630 ;
		LAYER M4 ;
		RECT 0.227 94.002 15.977 94.162 ;
		LAYER M4 ;
		RECT 0.227 94.910 15.977 95.070 ;
		LAYER M4 ;
		RECT 0.227 95.442 15.977 95.602 ;
		LAYER M4 ;
		RECT 0.227 96.350 15.977 96.510 ;
		LAYER M4 ;
		RECT 0.227 96.882 15.977 97.042 ;
		LAYER M4 ;
		RECT 0.227 97.790 15.977 97.950 ;
		LAYER M4 ;
		RECT 0.227 98.322 15.977 98.482 ;
		LAYER M4 ;
		RECT 0.227 99.230 15.977 99.390 ;
		LAYER M4 ;
		RECT 0.227 99.762 15.977 99.922 ;
		LAYER M4 ;
		RECT 0.227 100.670 15.977 100.830 ;
		LAYER M4 ;
		RECT 0.227 101.202 15.977 101.362 ;
		LAYER M4 ;
		RECT 0.227 102.110 15.977 102.270 ;
		LAYER M4 ;
		RECT 0.227 102.642 15.977 102.802 ;
		LAYER M4 ;
		RECT 0.227 103.550 15.977 103.710 ;
		LAYER M4 ;
		RECT 0.227 104.082 15.977 104.242 ;
		LAYER M4 ;
		RECT 0.227 104.990 15.977 105.150 ;
		LAYER M4 ;
		RECT 0.227 105.522 15.977 105.682 ;
		LAYER M4 ;
		RECT 0.227 106.430 15.977 106.590 ;
		LAYER M4 ;
		RECT 0.227 106.962 15.977 107.122 ;
		LAYER M4 ;
		RECT 0.227 107.870 15.977 108.030 ;
		LAYER M4 ;
		RECT 0.227 108.402 15.977 108.562 ;
		LAYER M4 ;
		RECT 0.227 109.310 15.977 109.470 ;
		LAYER M4 ;
		RECT 0.227 109.842 15.977 110.002 ;
		LAYER M4 ;
		RECT 0.227 110.750 15.977 110.910 ;
		LAYER M4 ;
		RECT 0.227 111.282 15.977 111.442 ;
		LAYER M4 ;
		RECT 0.227 112.076 16.407 112.276 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 16.957 112.800 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 16.957 112.800 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 16.957 112.800 ;
	END
END TS6N16FFCLLSVTA64X32M4FW

END LIBRARY
