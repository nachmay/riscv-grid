# Created by MC2 : Version 2013.12.00.f on 2025/06/18, 12:59:41

 
###############################################################################
#                                                    
#        Technology     : TSMC 16nm CMOS Logic FinFet (FFC) HKMG
#        Memory Type    : TSMC 16nm FFC Two Port Register File with d130 bit cell
#        Library Name   : ts6n16ffcllsvta16x32m2fw (user specify : ts6n16ffcllsvta16x32m2fw)
#        Library Version: 170a
#        Generated Time : 2025/06/18, 12:58:42
###############################################################################
# STATEMENT OF USE                                                             
#                                                                              
#  This information contains confidential and proprietary information of TSMC. 
# No part of this information may be reproduced, transmitted, transcribed,     
# stored in a retrieval system, or translated into any human or computer       
# language, in any form or by any means, electronic, mechanical, magnetic,     
# optical, chemical, manual, or otherwise, without the prior written permission
# of TSMC. This information was prepared for informational purpose and is for  
# use by TSMC's customers only. TSMC reserves the right to make changes in the 
# inforrmation at any time and without notice.                                 
###############################################################################
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
#                                                                              

MACRO TS6N16FFCLLSVTA16X32M2FW
	CLASS BLOCK ;
	FOREIGN TS6N16FFCLLSVTA16X32M2FW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 17.137 BY 66.720 ;
	SYMMETRY X Y ;
	PIN AA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 29.102 17.137 29.182 ;
			LAYER M2 ;
			RECT 16.889 29.102 17.137 29.182 ;
			LAYER M3 ;
			RECT 16.889 29.102 17.137 29.182 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[0]

	PIN AA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 32.294 17.137 32.374 ;
			LAYER M2 ;
			RECT 16.889 32.294 17.137 32.374 ;
			LAYER M3 ;
			RECT 16.889 32.294 17.137 32.374 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[1]

	PIN AA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 30.698 17.137 30.778 ;
			LAYER M2 ;
			RECT 16.889 30.698 17.137 30.778 ;
			LAYER M3 ;
			RECT 16.889 30.698 17.137 30.778 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[2]

	PIN AA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 32.066 17.137 32.146 ;
			LAYER M2 ;
			RECT 16.889 32.066 17.137 32.146 ;
			LAYER M3 ;
			RECT 16.889 32.066 17.137 32.146 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[3]

	PIN AB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 37.538 17.137 37.618 ;
			LAYER M2 ;
			RECT 16.889 37.538 17.137 37.618 ;
			LAYER M3 ;
			RECT 16.889 37.538 17.137 37.618 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[0]

	PIN AB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 34.346 17.137 34.426 ;
			LAYER M2 ;
			RECT 16.889 34.346 17.137 34.426 ;
			LAYER M3 ;
			RECT 16.889 34.346 17.137 34.426 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[1]

	PIN AB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 35.942 17.137 36.022 ;
			LAYER M2 ;
			RECT 16.889 35.942 17.137 36.022 ;
			LAYER M3 ;
			RECT 16.889 35.942 17.137 36.022 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[2]

	PIN AB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 34.574 17.137 34.654 ;
			LAYER M2 ;
			RECT 16.889 34.574 17.137 34.654 ;
			LAYER M3 ;
			RECT 16.889 34.574 17.137 34.654 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[3]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 1.088 17.137 1.168 ;
			LAYER M2 ;
			RECT 16.889 1.088 17.137 1.168 ;
			LAYER M3 ;
			RECT 16.889 1.088 17.137 1.168 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 2.528 17.137 2.608 ;
			LAYER M2 ;
			RECT 16.889 2.528 17.137 2.608 ;
			LAYER M3 ;
			RECT 16.889 2.528 17.137 2.608 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 3.968 17.137 4.048 ;
			LAYER M2 ;
			RECT 16.889 3.968 17.137 4.048 ;
			LAYER M3 ;
			RECT 16.889 3.968 17.137 4.048 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 5.408 17.137 5.488 ;
			LAYER M2 ;
			RECT 16.889 5.408 17.137 5.488 ;
			LAYER M3 ;
			RECT 16.889 5.408 17.137 5.488 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 6.848 17.137 6.928 ;
			LAYER M2 ;
			RECT 16.889 6.848 17.137 6.928 ;
			LAYER M3 ;
			RECT 16.889 6.848 17.137 6.928 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 8.288 17.137 8.368 ;
			LAYER M2 ;
			RECT 16.889 8.288 17.137 8.368 ;
			LAYER M3 ;
			RECT 16.889 8.288 17.137 8.368 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 9.728 17.137 9.808 ;
			LAYER M2 ;
			RECT 16.889 9.728 17.137 9.808 ;
			LAYER M3 ;
			RECT 16.889 9.728 17.137 9.808 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 11.168 17.137 11.248 ;
			LAYER M2 ;
			RECT 16.889 11.168 17.137 11.248 ;
			LAYER M3 ;
			RECT 16.889 11.168 17.137 11.248 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 12.608 17.137 12.688 ;
			LAYER M2 ;
			RECT 16.889 12.608 17.137 12.688 ;
			LAYER M3 ;
			RECT 16.889 12.608 17.137 12.688 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 14.048 17.137 14.128 ;
			LAYER M2 ;
			RECT 16.889 14.048 17.137 14.128 ;
			LAYER M3 ;
			RECT 16.889 14.048 17.137 14.128 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 15.488 17.137 15.568 ;
			LAYER M2 ;
			RECT 16.889 15.488 17.137 15.568 ;
			LAYER M3 ;
			RECT 16.889 15.488 17.137 15.568 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 16.928 17.137 17.008 ;
			LAYER M2 ;
			RECT 16.889 16.928 17.137 17.008 ;
			LAYER M3 ;
			RECT 16.889 16.928 17.137 17.008 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 18.368 17.137 18.448 ;
			LAYER M2 ;
			RECT 16.889 18.368 17.137 18.448 ;
			LAYER M3 ;
			RECT 16.889 18.368 17.137 18.448 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 19.808 17.137 19.888 ;
			LAYER M2 ;
			RECT 16.889 19.808 17.137 19.888 ;
			LAYER M3 ;
			RECT 16.889 19.808 17.137 19.888 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 21.248 17.137 21.328 ;
			LAYER M2 ;
			RECT 16.889 21.248 17.137 21.328 ;
			LAYER M3 ;
			RECT 16.889 21.248 17.137 21.328 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 22.688 17.137 22.768 ;
			LAYER M2 ;
			RECT 16.889 22.688 17.137 22.768 ;
			LAYER M3 ;
			RECT 16.889 22.688 17.137 22.768 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 43.952 17.137 44.032 ;
			LAYER M2 ;
			RECT 16.889 43.952 17.137 44.032 ;
			LAYER M3 ;
			RECT 16.889 43.952 17.137 44.032 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 45.392 17.137 45.472 ;
			LAYER M2 ;
			RECT 16.889 45.392 17.137 45.472 ;
			LAYER M3 ;
			RECT 16.889 45.392 17.137 45.472 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 46.832 17.137 46.912 ;
			LAYER M2 ;
			RECT 16.889 46.832 17.137 46.912 ;
			LAYER M3 ;
			RECT 16.889 46.832 17.137 46.912 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 48.272 17.137 48.352 ;
			LAYER M2 ;
			RECT 16.889 48.272 17.137 48.352 ;
			LAYER M3 ;
			RECT 16.889 48.272 17.137 48.352 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 49.712 17.137 49.792 ;
			LAYER M2 ;
			RECT 16.889 49.712 17.137 49.792 ;
			LAYER M3 ;
			RECT 16.889 49.712 17.137 49.792 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 51.152 17.137 51.232 ;
			LAYER M2 ;
			RECT 16.889 51.152 17.137 51.232 ;
			LAYER M3 ;
			RECT 16.889 51.152 17.137 51.232 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 52.592 17.137 52.672 ;
			LAYER M2 ;
			RECT 16.889 52.592 17.137 52.672 ;
			LAYER M3 ;
			RECT 16.889 52.592 17.137 52.672 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 54.032 17.137 54.112 ;
			LAYER M2 ;
			RECT 16.889 54.032 17.137 54.112 ;
			LAYER M3 ;
			RECT 16.889 54.032 17.137 54.112 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 55.472 17.137 55.552 ;
			LAYER M2 ;
			RECT 16.889 55.472 17.137 55.552 ;
			LAYER M3 ;
			RECT 16.889 55.472 17.137 55.552 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 56.912 17.137 56.992 ;
			LAYER M2 ;
			RECT 16.889 56.912 17.137 56.992 ;
			LAYER M3 ;
			RECT 16.889 56.912 17.137 56.992 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 58.352 17.137 58.432 ;
			LAYER M2 ;
			RECT 16.889 58.352 17.137 58.432 ;
			LAYER M3 ;
			RECT 16.889 58.352 17.137 58.432 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 59.792 17.137 59.872 ;
			LAYER M2 ;
			RECT 16.889 59.792 17.137 59.872 ;
			LAYER M3 ;
			RECT 16.889 59.792 17.137 59.872 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 61.232 17.137 61.312 ;
			LAYER M2 ;
			RECT 16.889 61.232 17.137 61.312 ;
			LAYER M3 ;
			RECT 16.889 61.232 17.137 61.312 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 62.672 17.137 62.752 ;
			LAYER M2 ;
			RECT 16.889 62.672 17.137 62.752 ;
			LAYER M3 ;
			RECT 16.889 62.672 17.137 62.752 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 64.112 17.137 64.192 ;
			LAYER M2 ;
			RECT 16.889 64.112 17.137 64.192 ;
			LAYER M3 ;
			RECT 16.889 64.112 17.137 64.192 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 65.552 17.137 65.632 ;
			LAYER M2 ;
			RECT 16.889 65.552 17.137 65.632 ;
			LAYER M3 ;
			RECT 16.889 65.552 17.137 65.632 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[31]

	PIN CLKR
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 40.274 17.137 40.354 ;
			LAYER M2 ;
			RECT 16.889 40.274 17.137 40.354 ;
			LAYER M3 ;
			RECT 16.889 40.274 17.137 40.354 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2280 LAYER M2 ;
		ANTENNAMAXAREACAR 40.1766 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0128 LAYER M3 ;
		ANTENNAMAXAREACAR 179.9160 LAYER M3 ;
	END CLKR

	PIN CLKW
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 25.682 17.137 25.762 ;
			LAYER M2 ;
			RECT 16.889 25.682 17.137 25.762 ;
			LAYER M3 ;
			RECT 16.889 25.682 17.137 25.762 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.4639 LAYER M2 ;
		ANTENNAMAXAREACAR 44.8112 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0082 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0159 LAYER M3 ;
		ANTENNAMAXAREACAR 150.9920 LAYER M3 ;
	END CLKW

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 2.240 17.137 2.320 ;
			LAYER M2 ;
			RECT 16.889 2.240 17.137 2.320 ;
			LAYER M3 ;
			RECT 16.889 2.240 17.137 2.320 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 3.680 17.137 3.760 ;
			LAYER M2 ;
			RECT 16.889 3.680 17.137 3.760 ;
			LAYER M3 ;
			RECT 16.889 3.680 17.137 3.760 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 5.120 17.137 5.200 ;
			LAYER M2 ;
			RECT 16.889 5.120 17.137 5.200 ;
			LAYER M3 ;
			RECT 16.889 5.120 17.137 5.200 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 6.560 17.137 6.640 ;
			LAYER M2 ;
			RECT 16.889 6.560 17.137 6.640 ;
			LAYER M3 ;
			RECT 16.889 6.560 17.137 6.640 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 8.000 17.137 8.080 ;
			LAYER M2 ;
			RECT 16.889 8.000 17.137 8.080 ;
			LAYER M3 ;
			RECT 16.889 8.000 17.137 8.080 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 9.440 17.137 9.520 ;
			LAYER M2 ;
			RECT 16.889 9.440 17.137 9.520 ;
			LAYER M3 ;
			RECT 16.889 9.440 17.137 9.520 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 10.880 17.137 10.960 ;
			LAYER M2 ;
			RECT 16.889 10.880 17.137 10.960 ;
			LAYER M3 ;
			RECT 16.889 10.880 17.137 10.960 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 12.320 17.137 12.400 ;
			LAYER M2 ;
			RECT 16.889 12.320 17.137 12.400 ;
			LAYER M3 ;
			RECT 16.889 12.320 17.137 12.400 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 13.760 17.137 13.840 ;
			LAYER M2 ;
			RECT 16.889 13.760 17.137 13.840 ;
			LAYER M3 ;
			RECT 16.889 13.760 17.137 13.840 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 15.200 17.137 15.280 ;
			LAYER M2 ;
			RECT 16.889 15.200 17.137 15.280 ;
			LAYER M3 ;
			RECT 16.889 15.200 17.137 15.280 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 16.640 17.137 16.720 ;
			LAYER M2 ;
			RECT 16.889 16.640 17.137 16.720 ;
			LAYER M3 ;
			RECT 16.889 16.640 17.137 16.720 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 18.080 17.137 18.160 ;
			LAYER M2 ;
			RECT 16.889 18.080 17.137 18.160 ;
			LAYER M3 ;
			RECT 16.889 18.080 17.137 18.160 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 19.520 17.137 19.600 ;
			LAYER M2 ;
			RECT 16.889 19.520 17.137 19.600 ;
			LAYER M3 ;
			RECT 16.889 19.520 17.137 19.600 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 20.960 17.137 21.040 ;
			LAYER M2 ;
			RECT 16.889 20.960 17.137 21.040 ;
			LAYER M3 ;
			RECT 16.889 20.960 17.137 21.040 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 22.400 17.137 22.480 ;
			LAYER M2 ;
			RECT 16.889 22.400 17.137 22.480 ;
			LAYER M3 ;
			RECT 16.889 22.400 17.137 22.480 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 23.840 17.137 23.920 ;
			LAYER M2 ;
			RECT 16.889 23.840 17.137 23.920 ;
			LAYER M3 ;
			RECT 16.889 23.840 17.137 23.920 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 42.800 17.137 42.880 ;
			LAYER M2 ;
			RECT 16.889 42.800 17.137 42.880 ;
			LAYER M3 ;
			RECT 16.889 42.800 17.137 42.880 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 44.240 17.137 44.320 ;
			LAYER M2 ;
			RECT 16.889 44.240 17.137 44.320 ;
			LAYER M3 ;
			RECT 16.889 44.240 17.137 44.320 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 45.680 17.137 45.760 ;
			LAYER M2 ;
			RECT 16.889 45.680 17.137 45.760 ;
			LAYER M3 ;
			RECT 16.889 45.680 17.137 45.760 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 47.120 17.137 47.200 ;
			LAYER M2 ;
			RECT 16.889 47.120 17.137 47.200 ;
			LAYER M3 ;
			RECT 16.889 47.120 17.137 47.200 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 48.560 17.137 48.640 ;
			LAYER M2 ;
			RECT 16.889 48.560 17.137 48.640 ;
			LAYER M3 ;
			RECT 16.889 48.560 17.137 48.640 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 50.000 17.137 50.080 ;
			LAYER M2 ;
			RECT 16.889 50.000 17.137 50.080 ;
			LAYER M3 ;
			RECT 16.889 50.000 17.137 50.080 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 51.440 17.137 51.520 ;
			LAYER M2 ;
			RECT 16.889 51.440 17.137 51.520 ;
			LAYER M3 ;
			RECT 16.889 51.440 17.137 51.520 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 52.880 17.137 52.960 ;
			LAYER M2 ;
			RECT 16.889 52.880 17.137 52.960 ;
			LAYER M3 ;
			RECT 16.889 52.880 17.137 52.960 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 54.320 17.137 54.400 ;
			LAYER M2 ;
			RECT 16.889 54.320 17.137 54.400 ;
			LAYER M3 ;
			RECT 16.889 54.320 17.137 54.400 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 55.760 17.137 55.840 ;
			LAYER M2 ;
			RECT 16.889 55.760 17.137 55.840 ;
			LAYER M3 ;
			RECT 16.889 55.760 17.137 55.840 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 57.200 17.137 57.280 ;
			LAYER M2 ;
			RECT 16.889 57.200 17.137 57.280 ;
			LAYER M3 ;
			RECT 16.889 57.200 17.137 57.280 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 58.640 17.137 58.720 ;
			LAYER M2 ;
			RECT 16.889 58.640 17.137 58.720 ;
			LAYER M3 ;
			RECT 16.889 58.640 17.137 58.720 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 60.080 17.137 60.160 ;
			LAYER M2 ;
			RECT 16.889 60.080 17.137 60.160 ;
			LAYER M3 ;
			RECT 16.889 60.080 17.137 60.160 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 61.520 17.137 61.600 ;
			LAYER M2 ;
			RECT 16.889 61.520 17.137 61.600 ;
			LAYER M3 ;
			RECT 16.889 61.520 17.137 61.600 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 62.960 17.137 63.040 ;
			LAYER M2 ;
			RECT 16.889 62.960 17.137 63.040 ;
			LAYER M3 ;
			RECT 16.889 62.960 17.137 63.040 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 64.400 17.137 64.480 ;
			LAYER M2 ;
			RECT 16.889 64.400 17.137 64.480 ;
			LAYER M3 ;
			RECT 16.889 64.400 17.137 64.480 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[31]

	PIN KP[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 27.050 17.137 27.130 ;
			LAYER M2 ;
			RECT 16.889 27.050 17.137 27.130 ;
			LAYER M3 ;
			RECT 16.889 27.050 17.137 27.130 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[0]

	PIN KP[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 27.278 17.137 27.358 ;
			LAYER M2 ;
			RECT 16.889 27.278 17.137 27.358 ;
			LAYER M3 ;
			RECT 16.889 27.278 17.137 27.358 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[1]

	PIN KP[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 27.506 17.137 27.586 ;
			LAYER M2 ;
			RECT 16.889 27.506 17.137 27.586 ;
			LAYER M3 ;
			RECT 16.889 27.506 17.137 27.586 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[2]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 1.662 17.137 1.742 ;
			LAYER M2 ;
			RECT 16.889 1.662 17.137 1.742 ;
			LAYER M3 ;
			RECT 16.889 1.662 17.137 1.742 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 3.102 17.137 3.182 ;
			LAYER M2 ;
			RECT 16.889 3.102 17.137 3.182 ;
			LAYER M3 ;
			RECT 16.889 3.102 17.137 3.182 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 4.542 17.137 4.622 ;
			LAYER M2 ;
			RECT 16.889 4.542 17.137 4.622 ;
			LAYER M3 ;
			RECT 16.889 4.542 17.137 4.622 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 5.982 17.137 6.062 ;
			LAYER M2 ;
			RECT 16.889 5.982 17.137 6.062 ;
			LAYER M3 ;
			RECT 16.889 5.982 17.137 6.062 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 7.422 17.137 7.502 ;
			LAYER M2 ;
			RECT 16.889 7.422 17.137 7.502 ;
			LAYER M3 ;
			RECT 16.889 7.422 17.137 7.502 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 8.862 17.137 8.942 ;
			LAYER M2 ;
			RECT 16.889 8.862 17.137 8.942 ;
			LAYER M3 ;
			RECT 16.889 8.862 17.137 8.942 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 10.302 17.137 10.382 ;
			LAYER M2 ;
			RECT 16.889 10.302 17.137 10.382 ;
			LAYER M3 ;
			RECT 16.889 10.302 17.137 10.382 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 11.742 17.137 11.822 ;
			LAYER M2 ;
			RECT 16.889 11.742 17.137 11.822 ;
			LAYER M3 ;
			RECT 16.889 11.742 17.137 11.822 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 13.182 17.137 13.262 ;
			LAYER M2 ;
			RECT 16.889 13.182 17.137 13.262 ;
			LAYER M3 ;
			RECT 16.889 13.182 17.137 13.262 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 14.622 17.137 14.702 ;
			LAYER M2 ;
			RECT 16.889 14.622 17.137 14.702 ;
			LAYER M3 ;
			RECT 16.889 14.622 17.137 14.702 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 16.062 17.137 16.142 ;
			LAYER M2 ;
			RECT 16.889 16.062 17.137 16.142 ;
			LAYER M3 ;
			RECT 16.889 16.062 17.137 16.142 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 17.502 17.137 17.582 ;
			LAYER M2 ;
			RECT 16.889 17.502 17.137 17.582 ;
			LAYER M3 ;
			RECT 16.889 17.502 17.137 17.582 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 18.942 17.137 19.022 ;
			LAYER M2 ;
			RECT 16.889 18.942 17.137 19.022 ;
			LAYER M3 ;
			RECT 16.889 18.942 17.137 19.022 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 20.382 17.137 20.462 ;
			LAYER M2 ;
			RECT 16.889 20.382 17.137 20.462 ;
			LAYER M3 ;
			RECT 16.889 20.382 17.137 20.462 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 21.822 17.137 21.902 ;
			LAYER M2 ;
			RECT 16.889 21.822 17.137 21.902 ;
			LAYER M3 ;
			RECT 16.889 21.822 17.137 21.902 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 23.262 17.137 23.342 ;
			LAYER M2 ;
			RECT 16.889 23.262 17.137 23.342 ;
			LAYER M3 ;
			RECT 16.889 23.262 17.137 23.342 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 43.378 17.137 43.458 ;
			LAYER M2 ;
			RECT 16.889 43.378 17.137 43.458 ;
			LAYER M3 ;
			RECT 16.889 43.378 17.137 43.458 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 44.818 17.137 44.898 ;
			LAYER M2 ;
			RECT 16.889 44.818 17.137 44.898 ;
			LAYER M3 ;
			RECT 16.889 44.818 17.137 44.898 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 46.258 17.137 46.338 ;
			LAYER M2 ;
			RECT 16.889 46.258 17.137 46.338 ;
			LAYER M3 ;
			RECT 16.889 46.258 17.137 46.338 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 47.698 17.137 47.778 ;
			LAYER M2 ;
			RECT 16.889 47.698 17.137 47.778 ;
			LAYER M3 ;
			RECT 16.889 47.698 17.137 47.778 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 49.138 17.137 49.218 ;
			LAYER M2 ;
			RECT 16.889 49.138 17.137 49.218 ;
			LAYER M3 ;
			RECT 16.889 49.138 17.137 49.218 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 50.578 17.137 50.658 ;
			LAYER M2 ;
			RECT 16.889 50.578 17.137 50.658 ;
			LAYER M3 ;
			RECT 16.889 50.578 17.137 50.658 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 52.018 17.137 52.098 ;
			LAYER M2 ;
			RECT 16.889 52.018 17.137 52.098 ;
			LAYER M3 ;
			RECT 16.889 52.018 17.137 52.098 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 53.458 17.137 53.538 ;
			LAYER M2 ;
			RECT 16.889 53.458 17.137 53.538 ;
			LAYER M3 ;
			RECT 16.889 53.458 17.137 53.538 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 54.898 17.137 54.978 ;
			LAYER M2 ;
			RECT 16.889 54.898 17.137 54.978 ;
			LAYER M3 ;
			RECT 16.889 54.898 17.137 54.978 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 56.338 17.137 56.418 ;
			LAYER M2 ;
			RECT 16.889 56.338 17.137 56.418 ;
			LAYER M3 ;
			RECT 16.889 56.338 17.137 56.418 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 57.778 17.137 57.858 ;
			LAYER M2 ;
			RECT 16.889 57.778 17.137 57.858 ;
			LAYER M3 ;
			RECT 16.889 57.778 17.137 57.858 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 59.218 17.137 59.298 ;
			LAYER M2 ;
			RECT 16.889 59.218 17.137 59.298 ;
			LAYER M3 ;
			RECT 16.889 59.218 17.137 59.298 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 60.658 17.137 60.738 ;
			LAYER M2 ;
			RECT 16.889 60.658 17.137 60.738 ;
			LAYER M3 ;
			RECT 16.889 60.658 17.137 60.738 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 62.098 17.137 62.178 ;
			LAYER M2 ;
			RECT 16.889 62.098 17.137 62.178 ;
			LAYER M3 ;
			RECT 16.889 62.098 17.137 62.178 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 63.538 17.137 63.618 ;
			LAYER M2 ;
			RECT 16.889 63.538 17.137 63.618 ;
			LAYER M3 ;
			RECT 16.889 63.538 17.137 63.618 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 64.978 17.137 65.058 ;
			LAYER M2 ;
			RECT 16.889 64.978 17.137 65.058 ;
			LAYER M3 ;
			RECT 16.889 64.978 17.137 65.058 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[31]

	PIN RCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 42.098 17.137 42.178 ;
			LAYER M2 ;
			RECT 16.889 42.098 17.137 42.178 ;
			LAYER M3 ;
			RECT 16.889 42.098 17.137 42.178 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[0]

	PIN RCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 41.870 17.137 41.950 ;
			LAYER M2 ;
			RECT 16.889 41.870 17.137 41.950 ;
			LAYER M3 ;
			RECT 16.889 41.870 17.137 41.950 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[1]

	PIN REB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 38.450 17.137 38.530 ;
			LAYER M2 ;
			RECT 16.889 38.450 17.137 38.530 ;
			LAYER M3 ;
			RECT 16.889 38.450 17.137 38.530 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0860 LAYER M1 ;
		ANTENNAMAXAREACAR 12.8828 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0840 LAYER M2 ;
		ANTENNAMAXAREACAR 20.5069 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4602 LAYER M3 ;
		ANTENNAMAXAREACAR 218.8550 LAYER M3 ;
	END REB

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.624 17.017 1.784 ;
			LAYER M4 ;
			RECT 0.120 3.064 17.017 3.224 ;
			LAYER M4 ;
			RECT 0.120 4.504 17.017 4.664 ;
			LAYER M4 ;
			RECT 0.120 5.944 17.017 6.104 ;
			LAYER M4 ;
			RECT 0.120 7.384 17.017 7.544 ;
			LAYER M4 ;
			RECT 0.120 8.824 17.017 8.984 ;
			LAYER M4 ;
			RECT 0.120 10.264 17.017 10.424 ;
			LAYER M4 ;
			RECT 0.120 11.704 17.017 11.864 ;
			LAYER M4 ;
			RECT 0.120 13.144 17.017 13.304 ;
			LAYER M4 ;
			RECT 0.120 14.584 17.017 14.744 ;
			LAYER M4 ;
			RECT 0.120 16.024 17.017 16.184 ;
			LAYER M4 ;
			RECT 0.120 17.464 17.017 17.624 ;
			LAYER M4 ;
			RECT 0.120 18.904 17.017 19.064 ;
			LAYER M4 ;
			RECT 0.120 20.344 17.017 20.504 ;
			LAYER M4 ;
			RECT 0.120 21.784 17.017 21.944 ;
			LAYER M4 ;
			RECT 0.120 23.224 17.017 23.384 ;
			LAYER M4 ;
			RECT 0.120 24.644 17.017 24.844 ;
			LAYER M4 ;
			RECT 0.120 25.580 17.017 25.780 ;
			LAYER M4 ;
			RECT 0.120 27.116 17.017 27.316 ;
			LAYER M4 ;
			RECT 0.120 28.652 17.017 28.852 ;
			LAYER M4 ;
			RECT 0.120 30.188 17.017 30.388 ;
			LAYER M4 ;
			RECT 0.120 31.724 17.017 31.924 ;
			LAYER M4 ;
			RECT 0.120 33.260 17.017 33.460 ;
			LAYER M4 ;
			RECT 0.120 34.796 17.017 34.996 ;
			LAYER M4 ;
			RECT 0.120 36.332 17.017 36.532 ;
			LAYER M4 ;
			RECT 0.120 37.868 17.017 38.068 ;
			LAYER M4 ;
			RECT 0.120 39.404 17.017 39.604 ;
			LAYER M4 ;
			RECT 0.120 40.940 17.017 41.140 ;
			LAYER M4 ;
			RECT 0.120 41.876 17.017 42.076 ;
			LAYER M4 ;
			RECT 0.120 43.336 17.017 43.496 ;
			LAYER M4 ;
			RECT 0.120 44.776 17.017 44.936 ;
			LAYER M4 ;
			RECT 0.120 46.216 17.017 46.376 ;
			LAYER M4 ;
			RECT 0.120 47.656 17.017 47.816 ;
			LAYER M4 ;
			RECT 0.120 49.096 17.017 49.256 ;
			LAYER M4 ;
			RECT 0.120 50.536 17.017 50.696 ;
			LAYER M4 ;
			RECT 0.120 51.976 17.017 52.136 ;
			LAYER M4 ;
			RECT 0.120 53.416 17.017 53.576 ;
			LAYER M4 ;
			RECT 0.120 54.856 17.017 55.016 ;
			LAYER M4 ;
			RECT 0.120 56.296 17.017 56.456 ;
			LAYER M4 ;
			RECT 0.120 57.736 17.017 57.896 ;
			LAYER M4 ;
			RECT 0.120 59.176 17.017 59.336 ;
			LAYER M4 ;
			RECT 0.120 60.616 17.017 60.776 ;
			LAYER M4 ;
			RECT 0.120 62.056 17.017 62.216 ;
			LAYER M4 ;
			RECT 0.120 63.496 17.017 63.656 ;
			LAYER M4 ;
			RECT 0.120 64.936 17.017 65.096 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 0.884 17.017 1.084 ;
			LAYER M4 ;
			RECT 0.120 2.324 17.017 2.524 ;
			LAYER M4 ;
			RECT 0.120 3.764 17.017 3.964 ;
			LAYER M4 ;
			RECT 0.120 5.204 17.017 5.404 ;
			LAYER M4 ;
			RECT 0.120 6.644 17.017 6.844 ;
			LAYER M4 ;
			RECT 0.120 8.084 17.017 8.284 ;
			LAYER M4 ;
			RECT 0.120 9.524 17.017 9.724 ;
			LAYER M4 ;
			RECT 0.120 10.964 17.017 11.164 ;
			LAYER M4 ;
			RECT 0.120 12.404 17.017 12.604 ;
			LAYER M4 ;
			RECT 0.120 13.844 17.017 14.044 ;
			LAYER M4 ;
			RECT 0.120 15.284 17.017 15.484 ;
			LAYER M4 ;
			RECT 0.120 16.724 17.017 16.924 ;
			LAYER M4 ;
			RECT 0.120 18.164 17.017 18.364 ;
			LAYER M4 ;
			RECT 0.120 19.604 17.017 19.804 ;
			LAYER M4 ;
			RECT 0.120 21.044 17.017 21.244 ;
			LAYER M4 ;
			RECT 0.120 22.484 17.017 22.684 ;
			LAYER M4 ;
			RECT 0.120 23.924 17.017 24.124 ;
			LAYER M4 ;
			RECT 0.120 26.348 17.017 26.548 ;
			LAYER M4 ;
			RECT 0.120 27.884 17.017 28.084 ;
			LAYER M4 ;
			RECT 0.120 29.420 17.017 29.620 ;
			LAYER M4 ;
			RECT 0.120 30.956 17.017 31.156 ;
			LAYER M4 ;
			RECT 0.120 32.492 17.017 32.692 ;
			LAYER M4 ;
			RECT 0.120 34.028 17.017 34.228 ;
			LAYER M4 ;
			RECT 0.120 35.564 17.017 35.764 ;
			LAYER M4 ;
			RECT 0.120 37.100 17.017 37.300 ;
			LAYER M4 ;
			RECT 0.120 38.636 17.017 38.836 ;
			LAYER M4 ;
			RECT 0.120 40.172 17.017 40.372 ;
			LAYER M4 ;
			RECT 0.120 42.596 17.017 42.796 ;
			LAYER M4 ;
			RECT 0.120 44.036 17.017 44.236 ;
			LAYER M4 ;
			RECT 0.120 45.476 17.017 45.676 ;
			LAYER M4 ;
			RECT 0.120 46.916 17.017 47.116 ;
			LAYER M4 ;
			RECT 0.120 48.356 17.017 48.556 ;
			LAYER M4 ;
			RECT 0.120 49.796 17.017 49.996 ;
			LAYER M4 ;
			RECT 0.120 51.236 17.017 51.436 ;
			LAYER M4 ;
			RECT 0.120 52.676 17.017 52.876 ;
			LAYER M4 ;
			RECT 0.120 54.116 17.017 54.316 ;
			LAYER M4 ;
			RECT 0.120 55.556 17.017 55.756 ;
			LAYER M4 ;
			RECT 0.120 56.996 17.017 57.196 ;
			LAYER M4 ;
			RECT 0.120 58.436 17.017 58.636 ;
			LAYER M4 ;
			RECT 0.120 59.876 17.017 60.076 ;
			LAYER M4 ;
			RECT 0.120 61.316 17.017 61.516 ;
			LAYER M4 ;
			RECT 0.120 62.756 17.017 62.956 ;
			LAYER M4 ;
			RECT 0.120 64.196 17.017 64.396 ;
			LAYER M4 ;
			RECT 0.120 65.636 17.017 65.836 ;
		END
	END VSS

	PIN WCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 24.998 17.137 25.078 ;
			LAYER M2 ;
			RECT 16.889 24.998 17.137 25.078 ;
			LAYER M3 ;
			RECT 16.889 24.998 17.137 25.078 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[0]

	PIN WCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 24.770 17.137 24.850 ;
			LAYER M2 ;
			RECT 16.889 24.770 17.137 24.850 ;
			LAYER M3 ;
			RECT 16.889 24.770 17.137 24.850 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.889 28.190 17.137 28.270 ;
			LAYER M2 ;
			RECT 16.889 28.190 17.137 28.270 ;
			LAYER M3 ;
			RECT 16.889 28.190 17.137 28.270 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0886 LAYER M1 ;
		ANTENNAMAXAREACAR 9.6368 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0833 LAYER M2 ;
		ANTENNAMAXAREACAR 13.2425 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4593 LAYER M3 ;
		ANTENNAMAXAREACAR 211.0720 LAYER M3 ;
	END WEB

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 17.137 66.720 ;
		LAYER M2 ;
		RECT 0.000 0.000 17.137 66.720 ;
		LAYER M3 ;
		RECT 0.000 0.000 17.137 66.720 ;
		LAYER M4 ;
		RECT 0.227 0.524 16.587 0.724 ;
		LAYER M4 ;
		RECT 0.227 1.358 16.157 1.518 ;
		LAYER M4 ;
		RECT 0.227 1.890 16.157 2.050 ;
		LAYER M4 ;
		RECT 0.227 2.798 16.157 2.958 ;
		LAYER M4 ;
		RECT 0.227 3.330 16.157 3.490 ;
		LAYER M4 ;
		RECT 0.227 4.238 16.157 4.398 ;
		LAYER M4 ;
		RECT 0.227 4.770 16.157 4.930 ;
		LAYER M4 ;
		RECT 0.227 5.678 16.157 5.838 ;
		LAYER M4 ;
		RECT 0.227 6.210 16.157 6.370 ;
		LAYER M4 ;
		RECT 0.227 7.118 16.157 7.278 ;
		LAYER M4 ;
		RECT 0.227 7.650 16.157 7.810 ;
		LAYER M4 ;
		RECT 0.227 8.558 16.157 8.718 ;
		LAYER M4 ;
		RECT 0.227 9.090 16.157 9.250 ;
		LAYER M4 ;
		RECT 0.227 9.998 16.157 10.158 ;
		LAYER M4 ;
		RECT 0.227 10.530 16.157 10.690 ;
		LAYER M4 ;
		RECT 0.227 11.438 16.157 11.598 ;
		LAYER M4 ;
		RECT 0.227 11.970 16.157 12.130 ;
		LAYER M4 ;
		RECT 0.227 12.878 16.157 13.038 ;
		LAYER M4 ;
		RECT 0.227 13.410 16.157 13.570 ;
		LAYER M4 ;
		RECT 0.227 14.318 16.157 14.478 ;
		LAYER M4 ;
		RECT 0.227 14.850 16.157 15.010 ;
		LAYER M4 ;
		RECT 0.227 15.758 16.157 15.918 ;
		LAYER M4 ;
		RECT 0.227 16.290 16.157 16.450 ;
		LAYER M4 ;
		RECT 0.227 17.198 16.157 17.358 ;
		LAYER M4 ;
		RECT 0.227 17.730 16.157 17.890 ;
		LAYER M4 ;
		RECT 0.227 18.638 16.157 18.798 ;
		LAYER M4 ;
		RECT 0.227 19.170 16.157 19.330 ;
		LAYER M4 ;
		RECT 0.227 20.078 16.157 20.238 ;
		LAYER M4 ;
		RECT 0.227 20.610 16.157 20.770 ;
		LAYER M4 ;
		RECT 0.227 21.518 16.157 21.678 ;
		LAYER M4 ;
		RECT 0.227 22.050 16.157 22.210 ;
		LAYER M4 ;
		RECT 0.227 22.958 16.157 23.118 ;
		LAYER M4 ;
		RECT 0.227 23.490 16.157 23.650 ;
		LAYER M4 ;
		RECT 0.227 24.284 16.157 24.484 ;
		LAYER M4 ;
		RECT 0.227 25.196 16.157 25.396 ;
		LAYER M4 ;
		RECT 0.227 25.964 16.157 26.164 ;
		LAYER M4 ;
		RECT 0.227 26.732 16.157 26.932 ;
		LAYER M4 ;
		RECT 0.227 27.500 16.157 27.700 ;
		LAYER M4 ;
		RECT 0.227 28.268 16.157 28.468 ;
		LAYER M4 ;
		RECT 0.227 29.036 16.157 29.236 ;
		LAYER M4 ;
		RECT 0.227 29.804 16.157 30.004 ;
		LAYER M4 ;
		RECT 0.227 30.572 16.157 30.772 ;
		LAYER M4 ;
		RECT 0.227 31.340 16.157 31.540 ;
		LAYER M4 ;
		RECT 0.227 32.108 16.157 32.308 ;
		LAYER M4 ;
		RECT 0.227 32.876 16.157 33.076 ;
		LAYER M4 ;
		RECT 0.227 33.644 16.157 33.844 ;
		LAYER M4 ;
		RECT 0.227 34.412 16.157 34.612 ;
		LAYER M4 ;
		RECT 0.227 35.180 16.157 35.380 ;
		LAYER M4 ;
		RECT 0.227 35.948 16.157 36.148 ;
		LAYER M4 ;
		RECT 0.227 36.716 16.157 36.916 ;
		LAYER M4 ;
		RECT 0.227 37.484 16.157 37.684 ;
		LAYER M4 ;
		RECT 0.227 38.252 16.157 38.452 ;
		LAYER M4 ;
		RECT 0.227 39.020 16.157 39.220 ;
		LAYER M4 ;
		RECT 0.227 39.788 16.157 39.988 ;
		LAYER M4 ;
		RECT 0.227 40.556 16.157 40.756 ;
		LAYER M4 ;
		RECT 0.227 41.324 16.157 41.524 ;
		LAYER M4 ;
		RECT 0.227 42.236 16.157 42.436 ;
		LAYER M4 ;
		RECT 0.227 43.070 16.157 43.230 ;
		LAYER M4 ;
		RECT 0.227 43.602 16.157 43.762 ;
		LAYER M4 ;
		RECT 0.227 44.510 16.157 44.670 ;
		LAYER M4 ;
		RECT 0.227 45.042 16.157 45.202 ;
		LAYER M4 ;
		RECT 0.227 45.950 16.157 46.110 ;
		LAYER M4 ;
		RECT 0.227 46.482 16.157 46.642 ;
		LAYER M4 ;
		RECT 0.227 47.390 16.157 47.550 ;
		LAYER M4 ;
		RECT 0.227 47.922 16.157 48.082 ;
		LAYER M4 ;
		RECT 0.227 48.830 16.157 48.990 ;
		LAYER M4 ;
		RECT 0.227 49.362 16.157 49.522 ;
		LAYER M4 ;
		RECT 0.227 50.270 16.157 50.430 ;
		LAYER M4 ;
		RECT 0.227 50.802 16.157 50.962 ;
		LAYER M4 ;
		RECT 0.227 51.710 16.157 51.870 ;
		LAYER M4 ;
		RECT 0.227 52.242 16.157 52.402 ;
		LAYER M4 ;
		RECT 0.227 53.150 16.157 53.310 ;
		LAYER M4 ;
		RECT 0.227 53.682 16.157 53.842 ;
		LAYER M4 ;
		RECT 0.227 54.590 16.157 54.750 ;
		LAYER M4 ;
		RECT 0.227 55.122 16.157 55.282 ;
		LAYER M4 ;
		RECT 0.227 56.030 16.157 56.190 ;
		LAYER M4 ;
		RECT 0.227 56.562 16.157 56.722 ;
		LAYER M4 ;
		RECT 0.227 57.470 16.157 57.630 ;
		LAYER M4 ;
		RECT 0.227 58.002 16.157 58.162 ;
		LAYER M4 ;
		RECT 0.227 58.910 16.157 59.070 ;
		LAYER M4 ;
		RECT 0.227 59.442 16.157 59.602 ;
		LAYER M4 ;
		RECT 0.227 60.350 16.157 60.510 ;
		LAYER M4 ;
		RECT 0.227 60.882 16.157 61.042 ;
		LAYER M4 ;
		RECT 0.227 61.790 16.157 61.950 ;
		LAYER M4 ;
		RECT 0.227 62.322 16.157 62.482 ;
		LAYER M4 ;
		RECT 0.227 63.230 16.157 63.390 ;
		LAYER M4 ;
		RECT 0.227 63.762 16.157 63.922 ;
		LAYER M4 ;
		RECT 0.227 64.670 16.157 64.830 ;
		LAYER M4 ;
		RECT 0.227 65.202 16.157 65.362 ;
		LAYER M4 ;
		RECT 0.227 65.996 16.587 66.196 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 17.137 66.720 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 17.137 66.720 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 17.137 66.720 ;
	END
END TS6N16FFCLLSVTA16X32M2FW

END LIBRARY
