# Created by MC2 : Version 2013.12.00.f on 2025/06/23, 09:41:45

#******************************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn16ffcll1prf_2013.12.00.120a 								*/
# Technology     : TSMC 16nm CMOS Logic FinFet Compact (FFC) HKMG                                                             */
# Memory Type    : TSMC 16nm FFC One Port Register File with d0907 bit cell                                        	     */
# Library Name   : ts5n16ffcllsvta8x128m1sw (user specify : TS5N16FFCLLSVTA8X128M1SW)				*/
# Library Version: 120a													*/
# Generated Time : 2025/06/23, 09:41:36										  	*/
#******************************************************************************************************************************/
#														    		*/
# STATEMENT OF USE												    		*/
#														    		*/
# This information contains confidential and proprietary information of TSMC.                                   		*/
# No part of this information may be reproduced, transmitted, transcribed,					     		*/
# stored in a retrieval system, or translated into any human or computer					    		*/
# language, in any form or by any means, electronic, mechanical, magnetic,					    		*/
# optical, chemical, manual, or otherwise, without the prior written permission                                  		*/
# of TSMC. This information was prepared for informational purpose and is for				      			*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the				      		*/
# information at any time and without notice.								      			*/
#														 		*/
#******************************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS5N16FFCLLSVTA8X128M1SW
	CLASS BLOCK ;
	FOREIGN TS5N16FFCLLSVTA8X128M1SW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 16.009 BY 77.664 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 37.736 16.009 37.816 ;
			LAYER M2 ;
			RECT 15.761 37.736 16.009 37.816 ;
			LAYER M3 ;
			RECT 15.761 37.736 16.009 37.816 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.068400 LAYER M1 ;
		ANTENNAMAXAREACAR 3.793440 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.421680 LAYER M2 ;
		ANTENNAMAXAREACAR 21.112800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.772440 LAYER M3 ;
		ANTENNAMAXAREACAR 84.016600 LAYER M3 ;
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 37.160 16.009 37.240 ;
			LAYER M2 ;
			RECT 15.761 37.160 16.009 37.240 ;
			LAYER M3 ;
			RECT 15.761 37.160 16.009 37.240 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.068400 LAYER M1 ;
		ANTENNAMAXAREACAR 3.793440 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.421680 LAYER M2 ;
		ANTENNAMAXAREACAR 21.112800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.772440 LAYER M3 ;
		ANTENNAMAXAREACAR 84.016600 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 34.472 16.009 34.552 ;
			LAYER M2 ;
			RECT 15.761 34.472 16.009 34.552 ;
			LAYER M3 ;
			RECT 15.761 34.472 16.009 34.552 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.068400 LAYER M1 ;
		ANTENNAMAXAREACAR 3.793440 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.421680 LAYER M2 ;
		ANTENNAMAXAREACAR 21.112800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.772440 LAYER M3 ;
		ANTENNAMAXAREACAR 84.016600 LAYER M3 ;
	END A[2]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 1.356 16.009 1.436 ;
			LAYER M2 ;
			RECT 15.761 1.356 16.009 1.436 ;
			LAYER M3 ;
			RECT 15.761 1.356 16.009 1.436 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 1.540 16.009 1.620 ;
			LAYER M2 ;
			RECT 15.761 1.540 16.009 1.620 ;
			LAYER M3 ;
			RECT 15.761 1.540 16.009 1.620 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 2.364 16.009 2.444 ;
			LAYER M2 ;
			RECT 15.761 2.364 16.009 2.444 ;
			LAYER M3 ;
			RECT 15.761 2.364 16.009 2.444 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 2.548 16.009 2.628 ;
			LAYER M2 ;
			RECT 15.761 2.548 16.009 2.628 ;
			LAYER M3 ;
			RECT 15.761 2.548 16.009 2.628 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 3.372 16.009 3.452 ;
			LAYER M2 ;
			RECT 15.761 3.372 16.009 3.452 ;
			LAYER M3 ;
			RECT 15.761 3.372 16.009 3.452 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 3.556 16.009 3.636 ;
			LAYER M2 ;
			RECT 15.761 3.556 16.009 3.636 ;
			LAYER M3 ;
			RECT 15.761 3.556 16.009 3.636 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 4.380 16.009 4.460 ;
			LAYER M2 ;
			RECT 15.761 4.380 16.009 4.460 ;
			LAYER M3 ;
			RECT 15.761 4.380 16.009 4.460 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 4.564 16.009 4.644 ;
			LAYER M2 ;
			RECT 15.761 4.564 16.009 4.644 ;
			LAYER M3 ;
			RECT 15.761 4.564 16.009 4.644 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 5.388 16.009 5.468 ;
			LAYER M2 ;
			RECT 15.761 5.388 16.009 5.468 ;
			LAYER M3 ;
			RECT 15.761 5.388 16.009 5.468 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 5.572 16.009 5.652 ;
			LAYER M2 ;
			RECT 15.761 5.572 16.009 5.652 ;
			LAYER M3 ;
			RECT 15.761 5.572 16.009 5.652 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 6.396 16.009 6.476 ;
			LAYER M2 ;
			RECT 15.761 6.396 16.009 6.476 ;
			LAYER M3 ;
			RECT 15.761 6.396 16.009 6.476 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 6.580 16.009 6.660 ;
			LAYER M2 ;
			RECT 15.761 6.580 16.009 6.660 ;
			LAYER M3 ;
			RECT 15.761 6.580 16.009 6.660 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 7.404 16.009 7.484 ;
			LAYER M2 ;
			RECT 15.761 7.404 16.009 7.484 ;
			LAYER M3 ;
			RECT 15.761 7.404 16.009 7.484 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 7.588 16.009 7.668 ;
			LAYER M2 ;
			RECT 15.761 7.588 16.009 7.668 ;
			LAYER M3 ;
			RECT 15.761 7.588 16.009 7.668 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 8.412 16.009 8.492 ;
			LAYER M2 ;
			RECT 15.761 8.412 16.009 8.492 ;
			LAYER M3 ;
			RECT 15.761 8.412 16.009 8.492 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 8.596 16.009 8.676 ;
			LAYER M2 ;
			RECT 15.761 8.596 16.009 8.676 ;
			LAYER M3 ;
			RECT 15.761 8.596 16.009 8.676 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 9.420 16.009 9.500 ;
			LAYER M2 ;
			RECT 15.761 9.420 16.009 9.500 ;
			LAYER M3 ;
			RECT 15.761 9.420 16.009 9.500 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 9.604 16.009 9.684 ;
			LAYER M2 ;
			RECT 15.761 9.604 16.009 9.684 ;
			LAYER M3 ;
			RECT 15.761 9.604 16.009 9.684 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 10.428 16.009 10.508 ;
			LAYER M2 ;
			RECT 15.761 10.428 16.009 10.508 ;
			LAYER M3 ;
			RECT 15.761 10.428 16.009 10.508 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 10.612 16.009 10.692 ;
			LAYER M2 ;
			RECT 15.761 10.612 16.009 10.692 ;
			LAYER M3 ;
			RECT 15.761 10.612 16.009 10.692 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 11.436 16.009 11.516 ;
			LAYER M2 ;
			RECT 15.761 11.436 16.009 11.516 ;
			LAYER M3 ;
			RECT 15.761 11.436 16.009 11.516 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 11.620 16.009 11.700 ;
			LAYER M2 ;
			RECT 15.761 11.620 16.009 11.700 ;
			LAYER M3 ;
			RECT 15.761 11.620 16.009 11.700 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 12.444 16.009 12.524 ;
			LAYER M2 ;
			RECT 15.761 12.444 16.009 12.524 ;
			LAYER M3 ;
			RECT 15.761 12.444 16.009 12.524 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 12.628 16.009 12.708 ;
			LAYER M2 ;
			RECT 15.761 12.628 16.009 12.708 ;
			LAYER M3 ;
			RECT 15.761 12.628 16.009 12.708 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 13.452 16.009 13.532 ;
			LAYER M2 ;
			RECT 15.761 13.452 16.009 13.532 ;
			LAYER M3 ;
			RECT 15.761 13.452 16.009 13.532 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 13.636 16.009 13.716 ;
			LAYER M2 ;
			RECT 15.761 13.636 16.009 13.716 ;
			LAYER M3 ;
			RECT 15.761 13.636 16.009 13.716 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 14.460 16.009 14.540 ;
			LAYER M2 ;
			RECT 15.761 14.460 16.009 14.540 ;
			LAYER M3 ;
			RECT 15.761 14.460 16.009 14.540 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 14.644 16.009 14.724 ;
			LAYER M2 ;
			RECT 15.761 14.644 16.009 14.724 ;
			LAYER M3 ;
			RECT 15.761 14.644 16.009 14.724 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 15.468 16.009 15.548 ;
			LAYER M2 ;
			RECT 15.761 15.468 16.009 15.548 ;
			LAYER M3 ;
			RECT 15.761 15.468 16.009 15.548 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 15.652 16.009 15.732 ;
			LAYER M2 ;
			RECT 15.761 15.652 16.009 15.732 ;
			LAYER M3 ;
			RECT 15.761 15.652 16.009 15.732 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 16.476 16.009 16.556 ;
			LAYER M2 ;
			RECT 15.761 16.476 16.009 16.556 ;
			LAYER M3 ;
			RECT 15.761 16.476 16.009 16.556 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 16.660 16.009 16.740 ;
			LAYER M2 ;
			RECT 15.761 16.660 16.009 16.740 ;
			LAYER M3 ;
			RECT 15.761 16.660 16.009 16.740 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[31]

	PIN BWEB[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 17.484 16.009 17.564 ;
			LAYER M2 ;
			RECT 15.761 17.484 16.009 17.564 ;
			LAYER M3 ;
			RECT 15.761 17.484 16.009 17.564 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[32]

	PIN BWEB[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 17.668 16.009 17.748 ;
			LAYER M2 ;
			RECT 15.761 17.668 16.009 17.748 ;
			LAYER M3 ;
			RECT 15.761 17.668 16.009 17.748 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[33]

	PIN BWEB[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 18.492 16.009 18.572 ;
			LAYER M2 ;
			RECT 15.761 18.492 16.009 18.572 ;
			LAYER M3 ;
			RECT 15.761 18.492 16.009 18.572 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[34]

	PIN BWEB[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 18.676 16.009 18.756 ;
			LAYER M2 ;
			RECT 15.761 18.676 16.009 18.756 ;
			LAYER M3 ;
			RECT 15.761 18.676 16.009 18.756 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[35]

	PIN BWEB[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 19.500 16.009 19.580 ;
			LAYER M2 ;
			RECT 15.761 19.500 16.009 19.580 ;
			LAYER M3 ;
			RECT 15.761 19.500 16.009 19.580 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[36]

	PIN BWEB[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 19.684 16.009 19.764 ;
			LAYER M2 ;
			RECT 15.761 19.684 16.009 19.764 ;
			LAYER M3 ;
			RECT 15.761 19.684 16.009 19.764 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[37]

	PIN BWEB[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 20.508 16.009 20.588 ;
			LAYER M2 ;
			RECT 15.761 20.508 16.009 20.588 ;
			LAYER M3 ;
			RECT 15.761 20.508 16.009 20.588 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[38]

	PIN BWEB[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 20.692 16.009 20.772 ;
			LAYER M2 ;
			RECT 15.761 20.692 16.009 20.772 ;
			LAYER M3 ;
			RECT 15.761 20.692 16.009 20.772 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[39]

	PIN BWEB[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 21.516 16.009 21.596 ;
			LAYER M2 ;
			RECT 15.761 21.516 16.009 21.596 ;
			LAYER M3 ;
			RECT 15.761 21.516 16.009 21.596 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[40]

	PIN BWEB[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 21.700 16.009 21.780 ;
			LAYER M2 ;
			RECT 15.761 21.700 16.009 21.780 ;
			LAYER M3 ;
			RECT 15.761 21.700 16.009 21.780 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[41]

	PIN BWEB[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 22.524 16.009 22.604 ;
			LAYER M2 ;
			RECT 15.761 22.524 16.009 22.604 ;
			LAYER M3 ;
			RECT 15.761 22.524 16.009 22.604 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[42]

	PIN BWEB[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 22.708 16.009 22.788 ;
			LAYER M2 ;
			RECT 15.761 22.708 16.009 22.788 ;
			LAYER M3 ;
			RECT 15.761 22.708 16.009 22.788 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[43]

	PIN BWEB[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 23.532 16.009 23.612 ;
			LAYER M2 ;
			RECT 15.761 23.532 16.009 23.612 ;
			LAYER M3 ;
			RECT 15.761 23.532 16.009 23.612 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[44]

	PIN BWEB[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 23.716 16.009 23.796 ;
			LAYER M2 ;
			RECT 15.761 23.716 16.009 23.796 ;
			LAYER M3 ;
			RECT 15.761 23.716 16.009 23.796 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[45]

	PIN BWEB[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 24.540 16.009 24.620 ;
			LAYER M2 ;
			RECT 15.761 24.540 16.009 24.620 ;
			LAYER M3 ;
			RECT 15.761 24.540 16.009 24.620 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[46]

	PIN BWEB[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 24.724 16.009 24.804 ;
			LAYER M2 ;
			RECT 15.761 24.724 16.009 24.804 ;
			LAYER M3 ;
			RECT 15.761 24.724 16.009 24.804 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[47]

	PIN BWEB[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 25.548 16.009 25.628 ;
			LAYER M2 ;
			RECT 15.761 25.548 16.009 25.628 ;
			LAYER M3 ;
			RECT 15.761 25.548 16.009 25.628 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[48]

	PIN BWEB[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 25.732 16.009 25.812 ;
			LAYER M2 ;
			RECT 15.761 25.732 16.009 25.812 ;
			LAYER M3 ;
			RECT 15.761 25.732 16.009 25.812 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[49]

	PIN BWEB[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 26.556 16.009 26.636 ;
			LAYER M2 ;
			RECT 15.761 26.556 16.009 26.636 ;
			LAYER M3 ;
			RECT 15.761 26.556 16.009 26.636 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[50]

	PIN BWEB[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 26.740 16.009 26.820 ;
			LAYER M2 ;
			RECT 15.761 26.740 16.009 26.820 ;
			LAYER M3 ;
			RECT 15.761 26.740 16.009 26.820 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[51]

	PIN BWEB[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 27.564 16.009 27.644 ;
			LAYER M2 ;
			RECT 15.761 27.564 16.009 27.644 ;
			LAYER M3 ;
			RECT 15.761 27.564 16.009 27.644 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[52]

	PIN BWEB[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 27.748 16.009 27.828 ;
			LAYER M2 ;
			RECT 15.761 27.748 16.009 27.828 ;
			LAYER M3 ;
			RECT 15.761 27.748 16.009 27.828 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[53]

	PIN BWEB[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 28.572 16.009 28.652 ;
			LAYER M2 ;
			RECT 15.761 28.572 16.009 28.652 ;
			LAYER M3 ;
			RECT 15.761 28.572 16.009 28.652 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[54]

	PIN BWEB[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 28.756 16.009 28.836 ;
			LAYER M2 ;
			RECT 15.761 28.756 16.009 28.836 ;
			LAYER M3 ;
			RECT 15.761 28.756 16.009 28.836 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[55]

	PIN BWEB[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 29.580 16.009 29.660 ;
			LAYER M2 ;
			RECT 15.761 29.580 16.009 29.660 ;
			LAYER M3 ;
			RECT 15.761 29.580 16.009 29.660 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[56]

	PIN BWEB[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 29.764 16.009 29.844 ;
			LAYER M2 ;
			RECT 15.761 29.764 16.009 29.844 ;
			LAYER M3 ;
			RECT 15.761 29.764 16.009 29.844 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[57]

	PIN BWEB[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 30.588 16.009 30.668 ;
			LAYER M2 ;
			RECT 15.761 30.588 16.009 30.668 ;
			LAYER M3 ;
			RECT 15.761 30.588 16.009 30.668 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[58]

	PIN BWEB[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 30.772 16.009 30.852 ;
			LAYER M2 ;
			RECT 15.761 30.772 16.009 30.852 ;
			LAYER M3 ;
			RECT 15.761 30.772 16.009 30.852 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[59]

	PIN BWEB[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 31.596 16.009 31.676 ;
			LAYER M2 ;
			RECT 15.761 31.596 16.009 31.676 ;
			LAYER M3 ;
			RECT 15.761 31.596 16.009 31.676 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[60]

	PIN BWEB[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 31.780 16.009 31.860 ;
			LAYER M2 ;
			RECT 15.761 31.780 16.009 31.860 ;
			LAYER M3 ;
			RECT 15.761 31.780 16.009 31.860 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[61]

	PIN BWEB[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 32.604 16.009 32.684 ;
			LAYER M2 ;
			RECT 15.761 32.604 16.009 32.684 ;
			LAYER M3 ;
			RECT 15.761 32.604 16.009 32.684 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[62]

	PIN BWEB[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 32.788 16.009 32.868 ;
			LAYER M2 ;
			RECT 15.761 32.788 16.009 32.868 ;
			LAYER M3 ;
			RECT 15.761 32.788 16.009 32.868 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[63]

	PIN BWEB[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 44.796 16.009 44.876 ;
			LAYER M2 ;
			RECT 15.761 44.796 16.009 44.876 ;
			LAYER M3 ;
			RECT 15.761 44.796 16.009 44.876 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[64]

	PIN BWEB[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 44.980 16.009 45.060 ;
			LAYER M2 ;
			RECT 15.761 44.980 16.009 45.060 ;
			LAYER M3 ;
			RECT 15.761 44.980 16.009 45.060 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[65]

	PIN BWEB[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 45.804 16.009 45.884 ;
			LAYER M2 ;
			RECT 15.761 45.804 16.009 45.884 ;
			LAYER M3 ;
			RECT 15.761 45.804 16.009 45.884 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[66]

	PIN BWEB[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 45.988 16.009 46.068 ;
			LAYER M2 ;
			RECT 15.761 45.988 16.009 46.068 ;
			LAYER M3 ;
			RECT 15.761 45.988 16.009 46.068 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[67]

	PIN BWEB[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 46.812 16.009 46.892 ;
			LAYER M2 ;
			RECT 15.761 46.812 16.009 46.892 ;
			LAYER M3 ;
			RECT 15.761 46.812 16.009 46.892 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[68]

	PIN BWEB[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 46.996 16.009 47.076 ;
			LAYER M2 ;
			RECT 15.761 46.996 16.009 47.076 ;
			LAYER M3 ;
			RECT 15.761 46.996 16.009 47.076 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[69]

	PIN BWEB[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 47.820 16.009 47.900 ;
			LAYER M2 ;
			RECT 15.761 47.820 16.009 47.900 ;
			LAYER M3 ;
			RECT 15.761 47.820 16.009 47.900 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[70]

	PIN BWEB[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 48.004 16.009 48.084 ;
			LAYER M2 ;
			RECT 15.761 48.004 16.009 48.084 ;
			LAYER M3 ;
			RECT 15.761 48.004 16.009 48.084 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[71]

	PIN BWEB[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 48.828 16.009 48.908 ;
			LAYER M2 ;
			RECT 15.761 48.828 16.009 48.908 ;
			LAYER M3 ;
			RECT 15.761 48.828 16.009 48.908 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[72]

	PIN BWEB[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 49.012 16.009 49.092 ;
			LAYER M2 ;
			RECT 15.761 49.012 16.009 49.092 ;
			LAYER M3 ;
			RECT 15.761 49.012 16.009 49.092 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[73]

	PIN BWEB[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 49.836 16.009 49.916 ;
			LAYER M2 ;
			RECT 15.761 49.836 16.009 49.916 ;
			LAYER M3 ;
			RECT 15.761 49.836 16.009 49.916 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[74]

	PIN BWEB[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 50.020 16.009 50.100 ;
			LAYER M2 ;
			RECT 15.761 50.020 16.009 50.100 ;
			LAYER M3 ;
			RECT 15.761 50.020 16.009 50.100 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[75]

	PIN BWEB[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 50.844 16.009 50.924 ;
			LAYER M2 ;
			RECT 15.761 50.844 16.009 50.924 ;
			LAYER M3 ;
			RECT 15.761 50.844 16.009 50.924 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[76]

	PIN BWEB[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 51.028 16.009 51.108 ;
			LAYER M2 ;
			RECT 15.761 51.028 16.009 51.108 ;
			LAYER M3 ;
			RECT 15.761 51.028 16.009 51.108 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[77]

	PIN BWEB[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 51.852 16.009 51.932 ;
			LAYER M2 ;
			RECT 15.761 51.852 16.009 51.932 ;
			LAYER M3 ;
			RECT 15.761 51.852 16.009 51.932 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[78]

	PIN BWEB[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 52.036 16.009 52.116 ;
			LAYER M2 ;
			RECT 15.761 52.036 16.009 52.116 ;
			LAYER M3 ;
			RECT 15.761 52.036 16.009 52.116 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[79]

	PIN BWEB[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 52.860 16.009 52.940 ;
			LAYER M2 ;
			RECT 15.761 52.860 16.009 52.940 ;
			LAYER M3 ;
			RECT 15.761 52.860 16.009 52.940 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[80]

	PIN BWEB[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 53.044 16.009 53.124 ;
			LAYER M2 ;
			RECT 15.761 53.044 16.009 53.124 ;
			LAYER M3 ;
			RECT 15.761 53.044 16.009 53.124 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[81]

	PIN BWEB[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 53.868 16.009 53.948 ;
			LAYER M2 ;
			RECT 15.761 53.868 16.009 53.948 ;
			LAYER M3 ;
			RECT 15.761 53.868 16.009 53.948 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[82]

	PIN BWEB[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 54.052 16.009 54.132 ;
			LAYER M2 ;
			RECT 15.761 54.052 16.009 54.132 ;
			LAYER M3 ;
			RECT 15.761 54.052 16.009 54.132 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[83]

	PIN BWEB[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 54.876 16.009 54.956 ;
			LAYER M2 ;
			RECT 15.761 54.876 16.009 54.956 ;
			LAYER M3 ;
			RECT 15.761 54.876 16.009 54.956 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[84]

	PIN BWEB[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 55.060 16.009 55.140 ;
			LAYER M2 ;
			RECT 15.761 55.060 16.009 55.140 ;
			LAYER M3 ;
			RECT 15.761 55.060 16.009 55.140 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[85]

	PIN BWEB[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 55.884 16.009 55.964 ;
			LAYER M2 ;
			RECT 15.761 55.884 16.009 55.964 ;
			LAYER M3 ;
			RECT 15.761 55.884 16.009 55.964 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[86]

	PIN BWEB[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 56.068 16.009 56.148 ;
			LAYER M2 ;
			RECT 15.761 56.068 16.009 56.148 ;
			LAYER M3 ;
			RECT 15.761 56.068 16.009 56.148 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[87]

	PIN BWEB[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 56.892 16.009 56.972 ;
			LAYER M2 ;
			RECT 15.761 56.892 16.009 56.972 ;
			LAYER M3 ;
			RECT 15.761 56.892 16.009 56.972 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[88]

	PIN BWEB[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 57.076 16.009 57.156 ;
			LAYER M2 ;
			RECT 15.761 57.076 16.009 57.156 ;
			LAYER M3 ;
			RECT 15.761 57.076 16.009 57.156 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[89]

	PIN BWEB[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 57.900 16.009 57.980 ;
			LAYER M2 ;
			RECT 15.761 57.900 16.009 57.980 ;
			LAYER M3 ;
			RECT 15.761 57.900 16.009 57.980 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[90]

	PIN BWEB[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 58.084 16.009 58.164 ;
			LAYER M2 ;
			RECT 15.761 58.084 16.009 58.164 ;
			LAYER M3 ;
			RECT 15.761 58.084 16.009 58.164 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[91]

	PIN BWEB[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 58.908 16.009 58.988 ;
			LAYER M2 ;
			RECT 15.761 58.908 16.009 58.988 ;
			LAYER M3 ;
			RECT 15.761 58.908 16.009 58.988 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[92]

	PIN BWEB[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 59.092 16.009 59.172 ;
			LAYER M2 ;
			RECT 15.761 59.092 16.009 59.172 ;
			LAYER M3 ;
			RECT 15.761 59.092 16.009 59.172 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[93]

	PIN BWEB[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 59.916 16.009 59.996 ;
			LAYER M2 ;
			RECT 15.761 59.916 16.009 59.996 ;
			LAYER M3 ;
			RECT 15.761 59.916 16.009 59.996 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[94]

	PIN BWEB[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 60.100 16.009 60.180 ;
			LAYER M2 ;
			RECT 15.761 60.100 16.009 60.180 ;
			LAYER M3 ;
			RECT 15.761 60.100 16.009 60.180 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[95]

	PIN BWEB[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 60.924 16.009 61.004 ;
			LAYER M2 ;
			RECT 15.761 60.924 16.009 61.004 ;
			LAYER M3 ;
			RECT 15.761 60.924 16.009 61.004 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[96]

	PIN BWEB[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 61.108 16.009 61.188 ;
			LAYER M2 ;
			RECT 15.761 61.108 16.009 61.188 ;
			LAYER M3 ;
			RECT 15.761 61.108 16.009 61.188 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[97]

	PIN BWEB[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 61.932 16.009 62.012 ;
			LAYER M2 ;
			RECT 15.761 61.932 16.009 62.012 ;
			LAYER M3 ;
			RECT 15.761 61.932 16.009 62.012 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[98]

	PIN BWEB[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 62.116 16.009 62.196 ;
			LAYER M2 ;
			RECT 15.761 62.116 16.009 62.196 ;
			LAYER M3 ;
			RECT 15.761 62.116 16.009 62.196 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[99]

	PIN BWEB[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 62.940 16.009 63.020 ;
			LAYER M2 ;
			RECT 15.761 62.940 16.009 63.020 ;
			LAYER M3 ;
			RECT 15.761 62.940 16.009 63.020 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[100]

	PIN BWEB[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 63.124 16.009 63.204 ;
			LAYER M2 ;
			RECT 15.761 63.124 16.009 63.204 ;
			LAYER M3 ;
			RECT 15.761 63.124 16.009 63.204 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[101]

	PIN BWEB[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 63.948 16.009 64.028 ;
			LAYER M2 ;
			RECT 15.761 63.948 16.009 64.028 ;
			LAYER M3 ;
			RECT 15.761 63.948 16.009 64.028 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[102]

	PIN BWEB[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 64.132 16.009 64.212 ;
			LAYER M2 ;
			RECT 15.761 64.132 16.009 64.212 ;
			LAYER M3 ;
			RECT 15.761 64.132 16.009 64.212 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[103]

	PIN BWEB[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 64.956 16.009 65.036 ;
			LAYER M2 ;
			RECT 15.761 64.956 16.009 65.036 ;
			LAYER M3 ;
			RECT 15.761 64.956 16.009 65.036 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[104]

	PIN BWEB[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 65.140 16.009 65.220 ;
			LAYER M2 ;
			RECT 15.761 65.140 16.009 65.220 ;
			LAYER M3 ;
			RECT 15.761 65.140 16.009 65.220 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[105]

	PIN BWEB[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 65.964 16.009 66.044 ;
			LAYER M2 ;
			RECT 15.761 65.964 16.009 66.044 ;
			LAYER M3 ;
			RECT 15.761 65.964 16.009 66.044 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[106]

	PIN BWEB[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 66.148 16.009 66.228 ;
			LAYER M2 ;
			RECT 15.761 66.148 16.009 66.228 ;
			LAYER M3 ;
			RECT 15.761 66.148 16.009 66.228 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[107]

	PIN BWEB[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 66.972 16.009 67.052 ;
			LAYER M2 ;
			RECT 15.761 66.972 16.009 67.052 ;
			LAYER M3 ;
			RECT 15.761 66.972 16.009 67.052 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[108]

	PIN BWEB[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 67.156 16.009 67.236 ;
			LAYER M2 ;
			RECT 15.761 67.156 16.009 67.236 ;
			LAYER M3 ;
			RECT 15.761 67.156 16.009 67.236 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[109]

	PIN BWEB[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 67.980 16.009 68.060 ;
			LAYER M2 ;
			RECT 15.761 67.980 16.009 68.060 ;
			LAYER M3 ;
			RECT 15.761 67.980 16.009 68.060 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[110]

	PIN BWEB[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 68.164 16.009 68.244 ;
			LAYER M2 ;
			RECT 15.761 68.164 16.009 68.244 ;
			LAYER M3 ;
			RECT 15.761 68.164 16.009 68.244 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[111]

	PIN BWEB[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 68.988 16.009 69.068 ;
			LAYER M2 ;
			RECT 15.761 68.988 16.009 69.068 ;
			LAYER M3 ;
			RECT 15.761 68.988 16.009 69.068 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[112]

	PIN BWEB[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 69.172 16.009 69.252 ;
			LAYER M2 ;
			RECT 15.761 69.172 16.009 69.252 ;
			LAYER M3 ;
			RECT 15.761 69.172 16.009 69.252 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[113]

	PIN BWEB[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 69.996 16.009 70.076 ;
			LAYER M2 ;
			RECT 15.761 69.996 16.009 70.076 ;
			LAYER M3 ;
			RECT 15.761 69.996 16.009 70.076 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[114]

	PIN BWEB[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 70.180 16.009 70.260 ;
			LAYER M2 ;
			RECT 15.761 70.180 16.009 70.260 ;
			LAYER M3 ;
			RECT 15.761 70.180 16.009 70.260 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[115]

	PIN BWEB[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 71.004 16.009 71.084 ;
			LAYER M2 ;
			RECT 15.761 71.004 16.009 71.084 ;
			LAYER M3 ;
			RECT 15.761 71.004 16.009 71.084 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[116]

	PIN BWEB[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 71.188 16.009 71.268 ;
			LAYER M2 ;
			RECT 15.761 71.188 16.009 71.268 ;
			LAYER M3 ;
			RECT 15.761 71.188 16.009 71.268 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[117]

	PIN BWEB[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 72.012 16.009 72.092 ;
			LAYER M2 ;
			RECT 15.761 72.012 16.009 72.092 ;
			LAYER M3 ;
			RECT 15.761 72.012 16.009 72.092 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[118]

	PIN BWEB[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 72.196 16.009 72.276 ;
			LAYER M2 ;
			RECT 15.761 72.196 16.009 72.276 ;
			LAYER M3 ;
			RECT 15.761 72.196 16.009 72.276 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[119]

	PIN BWEB[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 73.020 16.009 73.100 ;
			LAYER M2 ;
			RECT 15.761 73.020 16.009 73.100 ;
			LAYER M3 ;
			RECT 15.761 73.020 16.009 73.100 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[120]

	PIN BWEB[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 73.204 16.009 73.284 ;
			LAYER M2 ;
			RECT 15.761 73.204 16.009 73.284 ;
			LAYER M3 ;
			RECT 15.761 73.204 16.009 73.284 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[121]

	PIN BWEB[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 74.028 16.009 74.108 ;
			LAYER M2 ;
			RECT 15.761 74.028 16.009 74.108 ;
			LAYER M3 ;
			RECT 15.761 74.028 16.009 74.108 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[122]

	PIN BWEB[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 74.212 16.009 74.292 ;
			LAYER M2 ;
			RECT 15.761 74.212 16.009 74.292 ;
			LAYER M3 ;
			RECT 15.761 74.212 16.009 74.292 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[123]

	PIN BWEB[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 75.036 16.009 75.116 ;
			LAYER M2 ;
			RECT 15.761 75.036 16.009 75.116 ;
			LAYER M3 ;
			RECT 15.761 75.036 16.009 75.116 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[124]

	PIN BWEB[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 75.220 16.009 75.300 ;
			LAYER M2 ;
			RECT 15.761 75.220 16.009 75.300 ;
			LAYER M3 ;
			RECT 15.761 75.220 16.009 75.300 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[125]

	PIN BWEB[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 76.044 16.009 76.124 ;
			LAYER M2 ;
			RECT 15.761 76.044 16.009 76.124 ;
			LAYER M3 ;
			RECT 15.761 76.044 16.009 76.124 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[126]

	PIN BWEB[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 76.228 16.009 76.308 ;
			LAYER M2 ;
			RECT 15.761 76.228 16.009 76.308 ;
			LAYER M3 ;
			RECT 15.761 76.228 16.009 76.308 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.133680 LAYER M1 ;
		ANTENNAMAXAREACAR 12.295900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.786000 LAYER M2 ;
		ANTENNAMAXAREACAR 174.657000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.348480 LAYER M3 ;
		ANTENNAMAXAREACAR 230.817000 LAYER M3 ;
	END BWEB[127]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 38.120 16.009 38.200 ;
			LAYER M2 ;
			RECT 15.761 38.120 16.009 38.200 ;
			LAYER M3 ;
			RECT 15.761 38.120 16.009 38.200 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.075840 LAYER M1 ;
		ANTENNAMAXAREACAR 5.721480 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.302640 LAYER M2 ;
		ANTENNAMAXAREACAR 32.594800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.691080 LAYER M3 ;
		ANTENNAMAXAREACAR 195.580000 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 36.776 16.009 36.856 ;
			LAYER M2 ;
			RECT 15.761 36.776 16.009 36.856 ;
			LAYER M3 ;
			RECT 15.761 36.776 16.009 36.856 ;
		END
		ANTENNAGATEAREA 0.175917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.609600 LAYER M1 ;
		ANTENNAMAXAREACAR 3.871320 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.042960 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.362280 LAYER VIA1 ;
		ANTENNAGATEAREA 0.175917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 2.367120 LAYER M2 ;
		ANTENNAMAXAREACAR 70.244900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.027000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.652080 LAYER VIA2 ;
		ANTENNAGATEAREA 0.175917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.218200 LAYER M3 ;
		ANTENNAMAXAREACAR 79.541000 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 1.036 16.009 1.116 ;
			LAYER M2 ;
			RECT 15.761 1.036 16.009 1.116 ;
			LAYER M3 ;
			RECT 15.761 1.036 16.009 1.116 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 1.860 16.009 1.940 ;
			LAYER M2 ;
			RECT 15.761 1.860 16.009 1.940 ;
			LAYER M3 ;
			RECT 15.761 1.860 16.009 1.940 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 2.044 16.009 2.124 ;
			LAYER M2 ;
			RECT 15.761 2.044 16.009 2.124 ;
			LAYER M3 ;
			RECT 15.761 2.044 16.009 2.124 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 2.868 16.009 2.948 ;
			LAYER M2 ;
			RECT 15.761 2.868 16.009 2.948 ;
			LAYER M3 ;
			RECT 15.761 2.868 16.009 2.948 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 3.052 16.009 3.132 ;
			LAYER M2 ;
			RECT 15.761 3.052 16.009 3.132 ;
			LAYER M3 ;
			RECT 15.761 3.052 16.009 3.132 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 3.876 16.009 3.956 ;
			LAYER M2 ;
			RECT 15.761 3.876 16.009 3.956 ;
			LAYER M3 ;
			RECT 15.761 3.876 16.009 3.956 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 4.060 16.009 4.140 ;
			LAYER M2 ;
			RECT 15.761 4.060 16.009 4.140 ;
			LAYER M3 ;
			RECT 15.761 4.060 16.009 4.140 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 4.884 16.009 4.964 ;
			LAYER M2 ;
			RECT 15.761 4.884 16.009 4.964 ;
			LAYER M3 ;
			RECT 15.761 4.884 16.009 4.964 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 5.068 16.009 5.148 ;
			LAYER M2 ;
			RECT 15.761 5.068 16.009 5.148 ;
			LAYER M3 ;
			RECT 15.761 5.068 16.009 5.148 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 5.892 16.009 5.972 ;
			LAYER M2 ;
			RECT 15.761 5.892 16.009 5.972 ;
			LAYER M3 ;
			RECT 15.761 5.892 16.009 5.972 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 6.076 16.009 6.156 ;
			LAYER M2 ;
			RECT 15.761 6.076 16.009 6.156 ;
			LAYER M3 ;
			RECT 15.761 6.076 16.009 6.156 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 6.900 16.009 6.980 ;
			LAYER M2 ;
			RECT 15.761 6.900 16.009 6.980 ;
			LAYER M3 ;
			RECT 15.761 6.900 16.009 6.980 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 7.084 16.009 7.164 ;
			LAYER M2 ;
			RECT 15.761 7.084 16.009 7.164 ;
			LAYER M3 ;
			RECT 15.761 7.084 16.009 7.164 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 7.908 16.009 7.988 ;
			LAYER M2 ;
			RECT 15.761 7.908 16.009 7.988 ;
			LAYER M3 ;
			RECT 15.761 7.908 16.009 7.988 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 8.092 16.009 8.172 ;
			LAYER M2 ;
			RECT 15.761 8.092 16.009 8.172 ;
			LAYER M3 ;
			RECT 15.761 8.092 16.009 8.172 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 8.916 16.009 8.996 ;
			LAYER M2 ;
			RECT 15.761 8.916 16.009 8.996 ;
			LAYER M3 ;
			RECT 15.761 8.916 16.009 8.996 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 9.100 16.009 9.180 ;
			LAYER M2 ;
			RECT 15.761 9.100 16.009 9.180 ;
			LAYER M3 ;
			RECT 15.761 9.100 16.009 9.180 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 9.924 16.009 10.004 ;
			LAYER M2 ;
			RECT 15.761 9.924 16.009 10.004 ;
			LAYER M3 ;
			RECT 15.761 9.924 16.009 10.004 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 10.108 16.009 10.188 ;
			LAYER M2 ;
			RECT 15.761 10.108 16.009 10.188 ;
			LAYER M3 ;
			RECT 15.761 10.108 16.009 10.188 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 10.932 16.009 11.012 ;
			LAYER M2 ;
			RECT 15.761 10.932 16.009 11.012 ;
			LAYER M3 ;
			RECT 15.761 10.932 16.009 11.012 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 11.116 16.009 11.196 ;
			LAYER M2 ;
			RECT 15.761 11.116 16.009 11.196 ;
			LAYER M3 ;
			RECT 15.761 11.116 16.009 11.196 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 11.940 16.009 12.020 ;
			LAYER M2 ;
			RECT 15.761 11.940 16.009 12.020 ;
			LAYER M3 ;
			RECT 15.761 11.940 16.009 12.020 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 12.124 16.009 12.204 ;
			LAYER M2 ;
			RECT 15.761 12.124 16.009 12.204 ;
			LAYER M3 ;
			RECT 15.761 12.124 16.009 12.204 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 12.948 16.009 13.028 ;
			LAYER M2 ;
			RECT 15.761 12.948 16.009 13.028 ;
			LAYER M3 ;
			RECT 15.761 12.948 16.009 13.028 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 13.132 16.009 13.212 ;
			LAYER M2 ;
			RECT 15.761 13.132 16.009 13.212 ;
			LAYER M3 ;
			RECT 15.761 13.132 16.009 13.212 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 13.956 16.009 14.036 ;
			LAYER M2 ;
			RECT 15.761 13.956 16.009 14.036 ;
			LAYER M3 ;
			RECT 15.761 13.956 16.009 14.036 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 14.140 16.009 14.220 ;
			LAYER M2 ;
			RECT 15.761 14.140 16.009 14.220 ;
			LAYER M3 ;
			RECT 15.761 14.140 16.009 14.220 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 14.964 16.009 15.044 ;
			LAYER M2 ;
			RECT 15.761 14.964 16.009 15.044 ;
			LAYER M3 ;
			RECT 15.761 14.964 16.009 15.044 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 15.148 16.009 15.228 ;
			LAYER M2 ;
			RECT 15.761 15.148 16.009 15.228 ;
			LAYER M3 ;
			RECT 15.761 15.148 16.009 15.228 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 15.972 16.009 16.052 ;
			LAYER M2 ;
			RECT 15.761 15.972 16.009 16.052 ;
			LAYER M3 ;
			RECT 15.761 15.972 16.009 16.052 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 16.156 16.009 16.236 ;
			LAYER M2 ;
			RECT 15.761 16.156 16.009 16.236 ;
			LAYER M3 ;
			RECT 15.761 16.156 16.009 16.236 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 16.980 16.009 17.060 ;
			LAYER M2 ;
			RECT 15.761 16.980 16.009 17.060 ;
			LAYER M3 ;
			RECT 15.761 16.980 16.009 17.060 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 17.164 16.009 17.244 ;
			LAYER M2 ;
			RECT 15.761 17.164 16.009 17.244 ;
			LAYER M3 ;
			RECT 15.761 17.164 16.009 17.244 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 17.988 16.009 18.068 ;
			LAYER M2 ;
			RECT 15.761 17.988 16.009 18.068 ;
			LAYER M3 ;
			RECT 15.761 17.988 16.009 18.068 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 18.172 16.009 18.252 ;
			LAYER M2 ;
			RECT 15.761 18.172 16.009 18.252 ;
			LAYER M3 ;
			RECT 15.761 18.172 16.009 18.252 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 18.996 16.009 19.076 ;
			LAYER M2 ;
			RECT 15.761 18.996 16.009 19.076 ;
			LAYER M3 ;
			RECT 15.761 18.996 16.009 19.076 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[35]

	PIN D[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 19.180 16.009 19.260 ;
			LAYER M2 ;
			RECT 15.761 19.180 16.009 19.260 ;
			LAYER M3 ;
			RECT 15.761 19.180 16.009 19.260 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[36]

	PIN D[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 20.004 16.009 20.084 ;
			LAYER M2 ;
			RECT 15.761 20.004 16.009 20.084 ;
			LAYER M3 ;
			RECT 15.761 20.004 16.009 20.084 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[37]

	PIN D[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 20.188 16.009 20.268 ;
			LAYER M2 ;
			RECT 15.761 20.188 16.009 20.268 ;
			LAYER M3 ;
			RECT 15.761 20.188 16.009 20.268 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[38]

	PIN D[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 21.012 16.009 21.092 ;
			LAYER M2 ;
			RECT 15.761 21.012 16.009 21.092 ;
			LAYER M3 ;
			RECT 15.761 21.012 16.009 21.092 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[39]

	PIN D[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 21.196 16.009 21.276 ;
			LAYER M2 ;
			RECT 15.761 21.196 16.009 21.276 ;
			LAYER M3 ;
			RECT 15.761 21.196 16.009 21.276 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[40]

	PIN D[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 22.020 16.009 22.100 ;
			LAYER M2 ;
			RECT 15.761 22.020 16.009 22.100 ;
			LAYER M3 ;
			RECT 15.761 22.020 16.009 22.100 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[41]

	PIN D[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 22.204 16.009 22.284 ;
			LAYER M2 ;
			RECT 15.761 22.204 16.009 22.284 ;
			LAYER M3 ;
			RECT 15.761 22.204 16.009 22.284 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[42]

	PIN D[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 23.028 16.009 23.108 ;
			LAYER M2 ;
			RECT 15.761 23.028 16.009 23.108 ;
			LAYER M3 ;
			RECT 15.761 23.028 16.009 23.108 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[43]

	PIN D[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 23.212 16.009 23.292 ;
			LAYER M2 ;
			RECT 15.761 23.212 16.009 23.292 ;
			LAYER M3 ;
			RECT 15.761 23.212 16.009 23.292 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[44]

	PIN D[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 24.036 16.009 24.116 ;
			LAYER M2 ;
			RECT 15.761 24.036 16.009 24.116 ;
			LAYER M3 ;
			RECT 15.761 24.036 16.009 24.116 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[45]

	PIN D[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 24.220 16.009 24.300 ;
			LAYER M2 ;
			RECT 15.761 24.220 16.009 24.300 ;
			LAYER M3 ;
			RECT 15.761 24.220 16.009 24.300 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[46]

	PIN D[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 25.044 16.009 25.124 ;
			LAYER M2 ;
			RECT 15.761 25.044 16.009 25.124 ;
			LAYER M3 ;
			RECT 15.761 25.044 16.009 25.124 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[47]

	PIN D[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 25.228 16.009 25.308 ;
			LAYER M2 ;
			RECT 15.761 25.228 16.009 25.308 ;
			LAYER M3 ;
			RECT 15.761 25.228 16.009 25.308 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[48]

	PIN D[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 26.052 16.009 26.132 ;
			LAYER M2 ;
			RECT 15.761 26.052 16.009 26.132 ;
			LAYER M3 ;
			RECT 15.761 26.052 16.009 26.132 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[49]

	PIN D[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 26.236 16.009 26.316 ;
			LAYER M2 ;
			RECT 15.761 26.236 16.009 26.316 ;
			LAYER M3 ;
			RECT 15.761 26.236 16.009 26.316 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[50]

	PIN D[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 27.060 16.009 27.140 ;
			LAYER M2 ;
			RECT 15.761 27.060 16.009 27.140 ;
			LAYER M3 ;
			RECT 15.761 27.060 16.009 27.140 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[51]

	PIN D[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 27.244 16.009 27.324 ;
			LAYER M2 ;
			RECT 15.761 27.244 16.009 27.324 ;
			LAYER M3 ;
			RECT 15.761 27.244 16.009 27.324 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[52]

	PIN D[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 28.068 16.009 28.148 ;
			LAYER M2 ;
			RECT 15.761 28.068 16.009 28.148 ;
			LAYER M3 ;
			RECT 15.761 28.068 16.009 28.148 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[53]

	PIN D[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 28.252 16.009 28.332 ;
			LAYER M2 ;
			RECT 15.761 28.252 16.009 28.332 ;
			LAYER M3 ;
			RECT 15.761 28.252 16.009 28.332 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[54]

	PIN D[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 29.076 16.009 29.156 ;
			LAYER M2 ;
			RECT 15.761 29.076 16.009 29.156 ;
			LAYER M3 ;
			RECT 15.761 29.076 16.009 29.156 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[55]

	PIN D[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 29.260 16.009 29.340 ;
			LAYER M2 ;
			RECT 15.761 29.260 16.009 29.340 ;
			LAYER M3 ;
			RECT 15.761 29.260 16.009 29.340 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[56]

	PIN D[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 30.084 16.009 30.164 ;
			LAYER M2 ;
			RECT 15.761 30.084 16.009 30.164 ;
			LAYER M3 ;
			RECT 15.761 30.084 16.009 30.164 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[57]

	PIN D[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 30.268 16.009 30.348 ;
			LAYER M2 ;
			RECT 15.761 30.268 16.009 30.348 ;
			LAYER M3 ;
			RECT 15.761 30.268 16.009 30.348 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[58]

	PIN D[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 31.092 16.009 31.172 ;
			LAYER M2 ;
			RECT 15.761 31.092 16.009 31.172 ;
			LAYER M3 ;
			RECT 15.761 31.092 16.009 31.172 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[59]

	PIN D[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 31.276 16.009 31.356 ;
			LAYER M2 ;
			RECT 15.761 31.276 16.009 31.356 ;
			LAYER M3 ;
			RECT 15.761 31.276 16.009 31.356 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[60]

	PIN D[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 32.100 16.009 32.180 ;
			LAYER M2 ;
			RECT 15.761 32.100 16.009 32.180 ;
			LAYER M3 ;
			RECT 15.761 32.100 16.009 32.180 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[61]

	PIN D[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 32.284 16.009 32.364 ;
			LAYER M2 ;
			RECT 15.761 32.284 16.009 32.364 ;
			LAYER M3 ;
			RECT 15.761 32.284 16.009 32.364 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[62]

	PIN D[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 33.108 16.009 33.188 ;
			LAYER M2 ;
			RECT 15.761 33.108 16.009 33.188 ;
			LAYER M3 ;
			RECT 15.761 33.108 16.009 33.188 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[63]

	PIN D[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 44.476 16.009 44.556 ;
			LAYER M2 ;
			RECT 15.761 44.476 16.009 44.556 ;
			LAYER M3 ;
			RECT 15.761 44.476 16.009 44.556 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[64]

	PIN D[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 45.300 16.009 45.380 ;
			LAYER M2 ;
			RECT 15.761 45.300 16.009 45.380 ;
			LAYER M3 ;
			RECT 15.761 45.300 16.009 45.380 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[65]

	PIN D[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 45.484 16.009 45.564 ;
			LAYER M2 ;
			RECT 15.761 45.484 16.009 45.564 ;
			LAYER M3 ;
			RECT 15.761 45.484 16.009 45.564 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[66]

	PIN D[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 46.308 16.009 46.388 ;
			LAYER M2 ;
			RECT 15.761 46.308 16.009 46.388 ;
			LAYER M3 ;
			RECT 15.761 46.308 16.009 46.388 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[67]

	PIN D[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 46.492 16.009 46.572 ;
			LAYER M2 ;
			RECT 15.761 46.492 16.009 46.572 ;
			LAYER M3 ;
			RECT 15.761 46.492 16.009 46.572 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[68]

	PIN D[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 47.316 16.009 47.396 ;
			LAYER M2 ;
			RECT 15.761 47.316 16.009 47.396 ;
			LAYER M3 ;
			RECT 15.761 47.316 16.009 47.396 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[69]

	PIN D[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 47.500 16.009 47.580 ;
			LAYER M2 ;
			RECT 15.761 47.500 16.009 47.580 ;
			LAYER M3 ;
			RECT 15.761 47.500 16.009 47.580 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[70]

	PIN D[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 48.324 16.009 48.404 ;
			LAYER M2 ;
			RECT 15.761 48.324 16.009 48.404 ;
			LAYER M3 ;
			RECT 15.761 48.324 16.009 48.404 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[71]

	PIN D[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 48.508 16.009 48.588 ;
			LAYER M2 ;
			RECT 15.761 48.508 16.009 48.588 ;
			LAYER M3 ;
			RECT 15.761 48.508 16.009 48.588 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[72]

	PIN D[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 49.332 16.009 49.412 ;
			LAYER M2 ;
			RECT 15.761 49.332 16.009 49.412 ;
			LAYER M3 ;
			RECT 15.761 49.332 16.009 49.412 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[73]

	PIN D[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 49.516 16.009 49.596 ;
			LAYER M2 ;
			RECT 15.761 49.516 16.009 49.596 ;
			LAYER M3 ;
			RECT 15.761 49.516 16.009 49.596 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[74]

	PIN D[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 50.340 16.009 50.420 ;
			LAYER M2 ;
			RECT 15.761 50.340 16.009 50.420 ;
			LAYER M3 ;
			RECT 15.761 50.340 16.009 50.420 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[75]

	PIN D[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 50.524 16.009 50.604 ;
			LAYER M2 ;
			RECT 15.761 50.524 16.009 50.604 ;
			LAYER M3 ;
			RECT 15.761 50.524 16.009 50.604 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[76]

	PIN D[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 51.348 16.009 51.428 ;
			LAYER M2 ;
			RECT 15.761 51.348 16.009 51.428 ;
			LAYER M3 ;
			RECT 15.761 51.348 16.009 51.428 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[77]

	PIN D[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 51.532 16.009 51.612 ;
			LAYER M2 ;
			RECT 15.761 51.532 16.009 51.612 ;
			LAYER M3 ;
			RECT 15.761 51.532 16.009 51.612 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[78]

	PIN D[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 52.356 16.009 52.436 ;
			LAYER M2 ;
			RECT 15.761 52.356 16.009 52.436 ;
			LAYER M3 ;
			RECT 15.761 52.356 16.009 52.436 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[79]

	PIN D[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 52.540 16.009 52.620 ;
			LAYER M2 ;
			RECT 15.761 52.540 16.009 52.620 ;
			LAYER M3 ;
			RECT 15.761 52.540 16.009 52.620 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[80]

	PIN D[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 53.364 16.009 53.444 ;
			LAYER M2 ;
			RECT 15.761 53.364 16.009 53.444 ;
			LAYER M3 ;
			RECT 15.761 53.364 16.009 53.444 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[81]

	PIN D[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 53.548 16.009 53.628 ;
			LAYER M2 ;
			RECT 15.761 53.548 16.009 53.628 ;
			LAYER M3 ;
			RECT 15.761 53.548 16.009 53.628 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[82]

	PIN D[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 54.372 16.009 54.452 ;
			LAYER M2 ;
			RECT 15.761 54.372 16.009 54.452 ;
			LAYER M3 ;
			RECT 15.761 54.372 16.009 54.452 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[83]

	PIN D[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 54.556 16.009 54.636 ;
			LAYER M2 ;
			RECT 15.761 54.556 16.009 54.636 ;
			LAYER M3 ;
			RECT 15.761 54.556 16.009 54.636 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[84]

	PIN D[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 55.380 16.009 55.460 ;
			LAYER M2 ;
			RECT 15.761 55.380 16.009 55.460 ;
			LAYER M3 ;
			RECT 15.761 55.380 16.009 55.460 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[85]

	PIN D[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 55.564 16.009 55.644 ;
			LAYER M2 ;
			RECT 15.761 55.564 16.009 55.644 ;
			LAYER M3 ;
			RECT 15.761 55.564 16.009 55.644 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[86]

	PIN D[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 56.388 16.009 56.468 ;
			LAYER M2 ;
			RECT 15.761 56.388 16.009 56.468 ;
			LAYER M3 ;
			RECT 15.761 56.388 16.009 56.468 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[87]

	PIN D[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 56.572 16.009 56.652 ;
			LAYER M2 ;
			RECT 15.761 56.572 16.009 56.652 ;
			LAYER M3 ;
			RECT 15.761 56.572 16.009 56.652 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[88]

	PIN D[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 57.396 16.009 57.476 ;
			LAYER M2 ;
			RECT 15.761 57.396 16.009 57.476 ;
			LAYER M3 ;
			RECT 15.761 57.396 16.009 57.476 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[89]

	PIN D[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 57.580 16.009 57.660 ;
			LAYER M2 ;
			RECT 15.761 57.580 16.009 57.660 ;
			LAYER M3 ;
			RECT 15.761 57.580 16.009 57.660 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[90]

	PIN D[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 58.404 16.009 58.484 ;
			LAYER M2 ;
			RECT 15.761 58.404 16.009 58.484 ;
			LAYER M3 ;
			RECT 15.761 58.404 16.009 58.484 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[91]

	PIN D[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 58.588 16.009 58.668 ;
			LAYER M2 ;
			RECT 15.761 58.588 16.009 58.668 ;
			LAYER M3 ;
			RECT 15.761 58.588 16.009 58.668 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[92]

	PIN D[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 59.412 16.009 59.492 ;
			LAYER M2 ;
			RECT 15.761 59.412 16.009 59.492 ;
			LAYER M3 ;
			RECT 15.761 59.412 16.009 59.492 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[93]

	PIN D[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 59.596 16.009 59.676 ;
			LAYER M2 ;
			RECT 15.761 59.596 16.009 59.676 ;
			LAYER M3 ;
			RECT 15.761 59.596 16.009 59.676 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[94]

	PIN D[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 60.420 16.009 60.500 ;
			LAYER M2 ;
			RECT 15.761 60.420 16.009 60.500 ;
			LAYER M3 ;
			RECT 15.761 60.420 16.009 60.500 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[95]

	PIN D[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 60.604 16.009 60.684 ;
			LAYER M2 ;
			RECT 15.761 60.604 16.009 60.684 ;
			LAYER M3 ;
			RECT 15.761 60.604 16.009 60.684 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[96]

	PIN D[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 61.428 16.009 61.508 ;
			LAYER M2 ;
			RECT 15.761 61.428 16.009 61.508 ;
			LAYER M3 ;
			RECT 15.761 61.428 16.009 61.508 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[97]

	PIN D[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 61.612 16.009 61.692 ;
			LAYER M2 ;
			RECT 15.761 61.612 16.009 61.692 ;
			LAYER M3 ;
			RECT 15.761 61.612 16.009 61.692 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[98]

	PIN D[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 62.436 16.009 62.516 ;
			LAYER M2 ;
			RECT 15.761 62.436 16.009 62.516 ;
			LAYER M3 ;
			RECT 15.761 62.436 16.009 62.516 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[99]

	PIN D[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 62.620 16.009 62.700 ;
			LAYER M2 ;
			RECT 15.761 62.620 16.009 62.700 ;
			LAYER M3 ;
			RECT 15.761 62.620 16.009 62.700 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[100]

	PIN D[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 63.444 16.009 63.524 ;
			LAYER M2 ;
			RECT 15.761 63.444 16.009 63.524 ;
			LAYER M3 ;
			RECT 15.761 63.444 16.009 63.524 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[101]

	PIN D[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 63.628 16.009 63.708 ;
			LAYER M2 ;
			RECT 15.761 63.628 16.009 63.708 ;
			LAYER M3 ;
			RECT 15.761 63.628 16.009 63.708 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[102]

	PIN D[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 64.452 16.009 64.532 ;
			LAYER M2 ;
			RECT 15.761 64.452 16.009 64.532 ;
			LAYER M3 ;
			RECT 15.761 64.452 16.009 64.532 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[103]

	PIN D[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 64.636 16.009 64.716 ;
			LAYER M2 ;
			RECT 15.761 64.636 16.009 64.716 ;
			LAYER M3 ;
			RECT 15.761 64.636 16.009 64.716 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[104]

	PIN D[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 65.460 16.009 65.540 ;
			LAYER M2 ;
			RECT 15.761 65.460 16.009 65.540 ;
			LAYER M3 ;
			RECT 15.761 65.460 16.009 65.540 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[105]

	PIN D[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 65.644 16.009 65.724 ;
			LAYER M2 ;
			RECT 15.761 65.644 16.009 65.724 ;
			LAYER M3 ;
			RECT 15.761 65.644 16.009 65.724 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[106]

	PIN D[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 66.468 16.009 66.548 ;
			LAYER M2 ;
			RECT 15.761 66.468 16.009 66.548 ;
			LAYER M3 ;
			RECT 15.761 66.468 16.009 66.548 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[107]

	PIN D[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 66.652 16.009 66.732 ;
			LAYER M2 ;
			RECT 15.761 66.652 16.009 66.732 ;
			LAYER M3 ;
			RECT 15.761 66.652 16.009 66.732 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[108]

	PIN D[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 67.476 16.009 67.556 ;
			LAYER M2 ;
			RECT 15.761 67.476 16.009 67.556 ;
			LAYER M3 ;
			RECT 15.761 67.476 16.009 67.556 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[109]

	PIN D[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 67.660 16.009 67.740 ;
			LAYER M2 ;
			RECT 15.761 67.660 16.009 67.740 ;
			LAYER M3 ;
			RECT 15.761 67.660 16.009 67.740 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[110]

	PIN D[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 68.484 16.009 68.564 ;
			LAYER M2 ;
			RECT 15.761 68.484 16.009 68.564 ;
			LAYER M3 ;
			RECT 15.761 68.484 16.009 68.564 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[111]

	PIN D[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 68.668 16.009 68.748 ;
			LAYER M2 ;
			RECT 15.761 68.668 16.009 68.748 ;
			LAYER M3 ;
			RECT 15.761 68.668 16.009 68.748 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[112]

	PIN D[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 69.492 16.009 69.572 ;
			LAYER M2 ;
			RECT 15.761 69.492 16.009 69.572 ;
			LAYER M3 ;
			RECT 15.761 69.492 16.009 69.572 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[113]

	PIN D[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 69.676 16.009 69.756 ;
			LAYER M2 ;
			RECT 15.761 69.676 16.009 69.756 ;
			LAYER M3 ;
			RECT 15.761 69.676 16.009 69.756 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[114]

	PIN D[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 70.500 16.009 70.580 ;
			LAYER M2 ;
			RECT 15.761 70.500 16.009 70.580 ;
			LAYER M3 ;
			RECT 15.761 70.500 16.009 70.580 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[115]

	PIN D[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 70.684 16.009 70.764 ;
			LAYER M2 ;
			RECT 15.761 70.684 16.009 70.764 ;
			LAYER M3 ;
			RECT 15.761 70.684 16.009 70.764 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[116]

	PIN D[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 71.508 16.009 71.588 ;
			LAYER M2 ;
			RECT 15.761 71.508 16.009 71.588 ;
			LAYER M3 ;
			RECT 15.761 71.508 16.009 71.588 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[117]

	PIN D[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 71.692 16.009 71.772 ;
			LAYER M2 ;
			RECT 15.761 71.692 16.009 71.772 ;
			LAYER M3 ;
			RECT 15.761 71.692 16.009 71.772 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[118]

	PIN D[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 72.516 16.009 72.596 ;
			LAYER M2 ;
			RECT 15.761 72.516 16.009 72.596 ;
			LAYER M3 ;
			RECT 15.761 72.516 16.009 72.596 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[119]

	PIN D[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 72.700 16.009 72.780 ;
			LAYER M2 ;
			RECT 15.761 72.700 16.009 72.780 ;
			LAYER M3 ;
			RECT 15.761 72.700 16.009 72.780 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[120]

	PIN D[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 73.524 16.009 73.604 ;
			LAYER M2 ;
			RECT 15.761 73.524 16.009 73.604 ;
			LAYER M3 ;
			RECT 15.761 73.524 16.009 73.604 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[121]

	PIN D[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 73.708 16.009 73.788 ;
			LAYER M2 ;
			RECT 15.761 73.708 16.009 73.788 ;
			LAYER M3 ;
			RECT 15.761 73.708 16.009 73.788 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[122]

	PIN D[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 74.532 16.009 74.612 ;
			LAYER M2 ;
			RECT 15.761 74.532 16.009 74.612 ;
			LAYER M3 ;
			RECT 15.761 74.532 16.009 74.612 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[123]

	PIN D[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 74.716 16.009 74.796 ;
			LAYER M2 ;
			RECT 15.761 74.716 16.009 74.796 ;
			LAYER M3 ;
			RECT 15.761 74.716 16.009 74.796 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[124]

	PIN D[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 75.540 16.009 75.620 ;
			LAYER M2 ;
			RECT 15.761 75.540 16.009 75.620 ;
			LAYER M3 ;
			RECT 15.761 75.540 16.009 75.620 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[125]

	PIN D[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 75.724 16.009 75.804 ;
			LAYER M2 ;
			RECT 15.761 75.724 16.009 75.804 ;
			LAYER M3 ;
			RECT 15.761 75.724 16.009 75.804 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[126]

	PIN D[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 76.548 16.009 76.628 ;
			LAYER M2 ;
			RECT 15.761 76.548 16.009 76.628 ;
			LAYER M3 ;
			RECT 15.761 76.548 16.009 76.628 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.159240 LAYER M1 ;
		ANTENNAMAXAREACAR 18.814100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.017160 LAYER VIA1 ;
		ANTENNAMAXAREACAR 2.118600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.824280 LAYER M2 ;
		ANTENNAMAXAREACAR 269.018000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA2 ;
		ANTENNAMAXAREACAR 3.707640 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.300960 LAYER M3 ;
		ANTENNAMAXAREACAR 312.384000 LAYER M3 ;
	END D[127]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 1.196 16.009 1.276 ;
			LAYER M2 ;
			RECT 15.761 1.196 16.009 1.276 ;
			LAYER M3 ;
			RECT 15.761 1.196 16.009 1.276 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 1.700 16.009 1.780 ;
			LAYER M2 ;
			RECT 15.761 1.700 16.009 1.780 ;
			LAYER M3 ;
			RECT 15.761 1.700 16.009 1.780 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 2.204 16.009 2.284 ;
			LAYER M2 ;
			RECT 15.761 2.204 16.009 2.284 ;
			LAYER M3 ;
			RECT 15.761 2.204 16.009 2.284 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 2.708 16.009 2.788 ;
			LAYER M2 ;
			RECT 15.761 2.708 16.009 2.788 ;
			LAYER M3 ;
			RECT 15.761 2.708 16.009 2.788 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 3.212 16.009 3.292 ;
			LAYER M2 ;
			RECT 15.761 3.212 16.009 3.292 ;
			LAYER M3 ;
			RECT 15.761 3.212 16.009 3.292 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 3.716 16.009 3.796 ;
			LAYER M2 ;
			RECT 15.761 3.716 16.009 3.796 ;
			LAYER M3 ;
			RECT 15.761 3.716 16.009 3.796 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 4.220 16.009 4.300 ;
			LAYER M2 ;
			RECT 15.761 4.220 16.009 4.300 ;
			LAYER M3 ;
			RECT 15.761 4.220 16.009 4.300 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 4.724 16.009 4.804 ;
			LAYER M2 ;
			RECT 15.761 4.724 16.009 4.804 ;
			LAYER M3 ;
			RECT 15.761 4.724 16.009 4.804 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 5.228 16.009 5.308 ;
			LAYER M2 ;
			RECT 15.761 5.228 16.009 5.308 ;
			LAYER M3 ;
			RECT 15.761 5.228 16.009 5.308 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 5.732 16.009 5.812 ;
			LAYER M2 ;
			RECT 15.761 5.732 16.009 5.812 ;
			LAYER M3 ;
			RECT 15.761 5.732 16.009 5.812 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 6.236 16.009 6.316 ;
			LAYER M2 ;
			RECT 15.761 6.236 16.009 6.316 ;
			LAYER M3 ;
			RECT 15.761 6.236 16.009 6.316 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 6.740 16.009 6.820 ;
			LAYER M2 ;
			RECT 15.761 6.740 16.009 6.820 ;
			LAYER M3 ;
			RECT 15.761 6.740 16.009 6.820 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 7.244 16.009 7.324 ;
			LAYER M2 ;
			RECT 15.761 7.244 16.009 7.324 ;
			LAYER M3 ;
			RECT 15.761 7.244 16.009 7.324 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 7.748 16.009 7.828 ;
			LAYER M2 ;
			RECT 15.761 7.748 16.009 7.828 ;
			LAYER M3 ;
			RECT 15.761 7.748 16.009 7.828 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 8.252 16.009 8.332 ;
			LAYER M2 ;
			RECT 15.761 8.252 16.009 8.332 ;
			LAYER M3 ;
			RECT 15.761 8.252 16.009 8.332 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 8.756 16.009 8.836 ;
			LAYER M2 ;
			RECT 15.761 8.756 16.009 8.836 ;
			LAYER M3 ;
			RECT 15.761 8.756 16.009 8.836 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 9.260 16.009 9.340 ;
			LAYER M2 ;
			RECT 15.761 9.260 16.009 9.340 ;
			LAYER M3 ;
			RECT 15.761 9.260 16.009 9.340 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 9.764 16.009 9.844 ;
			LAYER M2 ;
			RECT 15.761 9.764 16.009 9.844 ;
			LAYER M3 ;
			RECT 15.761 9.764 16.009 9.844 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 10.268 16.009 10.348 ;
			LAYER M2 ;
			RECT 15.761 10.268 16.009 10.348 ;
			LAYER M3 ;
			RECT 15.761 10.268 16.009 10.348 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 10.772 16.009 10.852 ;
			LAYER M2 ;
			RECT 15.761 10.772 16.009 10.852 ;
			LAYER M3 ;
			RECT 15.761 10.772 16.009 10.852 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 11.276 16.009 11.356 ;
			LAYER M2 ;
			RECT 15.761 11.276 16.009 11.356 ;
			LAYER M3 ;
			RECT 15.761 11.276 16.009 11.356 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 11.780 16.009 11.860 ;
			LAYER M2 ;
			RECT 15.761 11.780 16.009 11.860 ;
			LAYER M3 ;
			RECT 15.761 11.780 16.009 11.860 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 12.284 16.009 12.364 ;
			LAYER M2 ;
			RECT 15.761 12.284 16.009 12.364 ;
			LAYER M3 ;
			RECT 15.761 12.284 16.009 12.364 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 12.788 16.009 12.868 ;
			LAYER M2 ;
			RECT 15.761 12.788 16.009 12.868 ;
			LAYER M3 ;
			RECT 15.761 12.788 16.009 12.868 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 13.292 16.009 13.372 ;
			LAYER M2 ;
			RECT 15.761 13.292 16.009 13.372 ;
			LAYER M3 ;
			RECT 15.761 13.292 16.009 13.372 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 13.796 16.009 13.876 ;
			LAYER M2 ;
			RECT 15.761 13.796 16.009 13.876 ;
			LAYER M3 ;
			RECT 15.761 13.796 16.009 13.876 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 14.300 16.009 14.380 ;
			LAYER M2 ;
			RECT 15.761 14.300 16.009 14.380 ;
			LAYER M3 ;
			RECT 15.761 14.300 16.009 14.380 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 14.804 16.009 14.884 ;
			LAYER M2 ;
			RECT 15.761 14.804 16.009 14.884 ;
			LAYER M3 ;
			RECT 15.761 14.804 16.009 14.884 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 15.308 16.009 15.388 ;
			LAYER M2 ;
			RECT 15.761 15.308 16.009 15.388 ;
			LAYER M3 ;
			RECT 15.761 15.308 16.009 15.388 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 15.812 16.009 15.892 ;
			LAYER M2 ;
			RECT 15.761 15.812 16.009 15.892 ;
			LAYER M3 ;
			RECT 15.761 15.812 16.009 15.892 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 16.316 16.009 16.396 ;
			LAYER M2 ;
			RECT 15.761 16.316 16.009 16.396 ;
			LAYER M3 ;
			RECT 15.761 16.316 16.009 16.396 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 16.820 16.009 16.900 ;
			LAYER M2 ;
			RECT 15.761 16.820 16.009 16.900 ;
			LAYER M3 ;
			RECT 15.761 16.820 16.009 16.900 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 17.324 16.009 17.404 ;
			LAYER M2 ;
			RECT 15.761 17.324 16.009 17.404 ;
			LAYER M3 ;
			RECT 15.761 17.324 16.009 17.404 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 17.828 16.009 17.908 ;
			LAYER M2 ;
			RECT 15.761 17.828 16.009 17.908 ;
			LAYER M3 ;
			RECT 15.761 17.828 16.009 17.908 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 18.332 16.009 18.412 ;
			LAYER M2 ;
			RECT 15.761 18.332 16.009 18.412 ;
			LAYER M3 ;
			RECT 15.761 18.332 16.009 18.412 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 18.836 16.009 18.916 ;
			LAYER M2 ;
			RECT 15.761 18.836 16.009 18.916 ;
			LAYER M3 ;
			RECT 15.761 18.836 16.009 18.916 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[35]

	PIN Q[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 19.340 16.009 19.420 ;
			LAYER M2 ;
			RECT 15.761 19.340 16.009 19.420 ;
			LAYER M3 ;
			RECT 15.761 19.340 16.009 19.420 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[36]

	PIN Q[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 19.844 16.009 19.924 ;
			LAYER M2 ;
			RECT 15.761 19.844 16.009 19.924 ;
			LAYER M3 ;
			RECT 15.761 19.844 16.009 19.924 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[37]

	PIN Q[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 20.348 16.009 20.428 ;
			LAYER M2 ;
			RECT 15.761 20.348 16.009 20.428 ;
			LAYER M3 ;
			RECT 15.761 20.348 16.009 20.428 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[38]

	PIN Q[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 20.852 16.009 20.932 ;
			LAYER M2 ;
			RECT 15.761 20.852 16.009 20.932 ;
			LAYER M3 ;
			RECT 15.761 20.852 16.009 20.932 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[39]

	PIN Q[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 21.356 16.009 21.436 ;
			LAYER M2 ;
			RECT 15.761 21.356 16.009 21.436 ;
			LAYER M3 ;
			RECT 15.761 21.356 16.009 21.436 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[40]

	PIN Q[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 21.860 16.009 21.940 ;
			LAYER M2 ;
			RECT 15.761 21.860 16.009 21.940 ;
			LAYER M3 ;
			RECT 15.761 21.860 16.009 21.940 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[41]

	PIN Q[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 22.364 16.009 22.444 ;
			LAYER M2 ;
			RECT 15.761 22.364 16.009 22.444 ;
			LAYER M3 ;
			RECT 15.761 22.364 16.009 22.444 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[42]

	PIN Q[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 22.868 16.009 22.948 ;
			LAYER M2 ;
			RECT 15.761 22.868 16.009 22.948 ;
			LAYER M3 ;
			RECT 15.761 22.868 16.009 22.948 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[43]

	PIN Q[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 23.372 16.009 23.452 ;
			LAYER M2 ;
			RECT 15.761 23.372 16.009 23.452 ;
			LAYER M3 ;
			RECT 15.761 23.372 16.009 23.452 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[44]

	PIN Q[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 23.876 16.009 23.956 ;
			LAYER M2 ;
			RECT 15.761 23.876 16.009 23.956 ;
			LAYER M3 ;
			RECT 15.761 23.876 16.009 23.956 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[45]

	PIN Q[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 24.380 16.009 24.460 ;
			LAYER M2 ;
			RECT 15.761 24.380 16.009 24.460 ;
			LAYER M3 ;
			RECT 15.761 24.380 16.009 24.460 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[46]

	PIN Q[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 24.884 16.009 24.964 ;
			LAYER M2 ;
			RECT 15.761 24.884 16.009 24.964 ;
			LAYER M3 ;
			RECT 15.761 24.884 16.009 24.964 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[47]

	PIN Q[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 25.388 16.009 25.468 ;
			LAYER M2 ;
			RECT 15.761 25.388 16.009 25.468 ;
			LAYER M3 ;
			RECT 15.761 25.388 16.009 25.468 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[48]

	PIN Q[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 25.892 16.009 25.972 ;
			LAYER M2 ;
			RECT 15.761 25.892 16.009 25.972 ;
			LAYER M3 ;
			RECT 15.761 25.892 16.009 25.972 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[49]

	PIN Q[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 26.396 16.009 26.476 ;
			LAYER M2 ;
			RECT 15.761 26.396 16.009 26.476 ;
			LAYER M3 ;
			RECT 15.761 26.396 16.009 26.476 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[50]

	PIN Q[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 26.900 16.009 26.980 ;
			LAYER M2 ;
			RECT 15.761 26.900 16.009 26.980 ;
			LAYER M3 ;
			RECT 15.761 26.900 16.009 26.980 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[51]

	PIN Q[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 27.404 16.009 27.484 ;
			LAYER M2 ;
			RECT 15.761 27.404 16.009 27.484 ;
			LAYER M3 ;
			RECT 15.761 27.404 16.009 27.484 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[52]

	PIN Q[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 27.908 16.009 27.988 ;
			LAYER M2 ;
			RECT 15.761 27.908 16.009 27.988 ;
			LAYER M3 ;
			RECT 15.761 27.908 16.009 27.988 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[53]

	PIN Q[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 28.412 16.009 28.492 ;
			LAYER M2 ;
			RECT 15.761 28.412 16.009 28.492 ;
			LAYER M3 ;
			RECT 15.761 28.412 16.009 28.492 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[54]

	PIN Q[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 28.916 16.009 28.996 ;
			LAYER M2 ;
			RECT 15.761 28.916 16.009 28.996 ;
			LAYER M3 ;
			RECT 15.761 28.916 16.009 28.996 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[55]

	PIN Q[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 29.420 16.009 29.500 ;
			LAYER M2 ;
			RECT 15.761 29.420 16.009 29.500 ;
			LAYER M3 ;
			RECT 15.761 29.420 16.009 29.500 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[56]

	PIN Q[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 29.924 16.009 30.004 ;
			LAYER M2 ;
			RECT 15.761 29.924 16.009 30.004 ;
			LAYER M3 ;
			RECT 15.761 29.924 16.009 30.004 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[57]

	PIN Q[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 30.428 16.009 30.508 ;
			LAYER M2 ;
			RECT 15.761 30.428 16.009 30.508 ;
			LAYER M3 ;
			RECT 15.761 30.428 16.009 30.508 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[58]

	PIN Q[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 30.932 16.009 31.012 ;
			LAYER M2 ;
			RECT 15.761 30.932 16.009 31.012 ;
			LAYER M3 ;
			RECT 15.761 30.932 16.009 31.012 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[59]

	PIN Q[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 31.436 16.009 31.516 ;
			LAYER M2 ;
			RECT 15.761 31.436 16.009 31.516 ;
			LAYER M3 ;
			RECT 15.761 31.436 16.009 31.516 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[60]

	PIN Q[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 31.940 16.009 32.020 ;
			LAYER M2 ;
			RECT 15.761 31.940 16.009 32.020 ;
			LAYER M3 ;
			RECT 15.761 31.940 16.009 32.020 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[61]

	PIN Q[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 32.444 16.009 32.524 ;
			LAYER M2 ;
			RECT 15.761 32.444 16.009 32.524 ;
			LAYER M3 ;
			RECT 15.761 32.444 16.009 32.524 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[62]

	PIN Q[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 32.948 16.009 33.028 ;
			LAYER M2 ;
			RECT 15.761 32.948 16.009 33.028 ;
			LAYER M3 ;
			RECT 15.761 32.948 16.009 33.028 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[63]

	PIN Q[64]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 44.636 16.009 44.716 ;
			LAYER M2 ;
			RECT 15.761 44.636 16.009 44.716 ;
			LAYER M3 ;
			RECT 15.761 44.636 16.009 44.716 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[64]

	PIN Q[65]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 45.140 16.009 45.220 ;
			LAYER M2 ;
			RECT 15.761 45.140 16.009 45.220 ;
			LAYER M3 ;
			RECT 15.761 45.140 16.009 45.220 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[65]

	PIN Q[66]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 45.644 16.009 45.724 ;
			LAYER M2 ;
			RECT 15.761 45.644 16.009 45.724 ;
			LAYER M3 ;
			RECT 15.761 45.644 16.009 45.724 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[66]

	PIN Q[67]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 46.148 16.009 46.228 ;
			LAYER M2 ;
			RECT 15.761 46.148 16.009 46.228 ;
			LAYER M3 ;
			RECT 15.761 46.148 16.009 46.228 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[67]

	PIN Q[68]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 46.652 16.009 46.732 ;
			LAYER M2 ;
			RECT 15.761 46.652 16.009 46.732 ;
			LAYER M3 ;
			RECT 15.761 46.652 16.009 46.732 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[68]

	PIN Q[69]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 47.156 16.009 47.236 ;
			LAYER M2 ;
			RECT 15.761 47.156 16.009 47.236 ;
			LAYER M3 ;
			RECT 15.761 47.156 16.009 47.236 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[69]

	PIN Q[70]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 47.660 16.009 47.740 ;
			LAYER M2 ;
			RECT 15.761 47.660 16.009 47.740 ;
			LAYER M3 ;
			RECT 15.761 47.660 16.009 47.740 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[70]

	PIN Q[71]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 48.164 16.009 48.244 ;
			LAYER M2 ;
			RECT 15.761 48.164 16.009 48.244 ;
			LAYER M3 ;
			RECT 15.761 48.164 16.009 48.244 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[71]

	PIN Q[72]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 48.668 16.009 48.748 ;
			LAYER M2 ;
			RECT 15.761 48.668 16.009 48.748 ;
			LAYER M3 ;
			RECT 15.761 48.668 16.009 48.748 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[72]

	PIN Q[73]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 49.172 16.009 49.252 ;
			LAYER M2 ;
			RECT 15.761 49.172 16.009 49.252 ;
			LAYER M3 ;
			RECT 15.761 49.172 16.009 49.252 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[73]

	PIN Q[74]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 49.676 16.009 49.756 ;
			LAYER M2 ;
			RECT 15.761 49.676 16.009 49.756 ;
			LAYER M3 ;
			RECT 15.761 49.676 16.009 49.756 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[74]

	PIN Q[75]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 50.180 16.009 50.260 ;
			LAYER M2 ;
			RECT 15.761 50.180 16.009 50.260 ;
			LAYER M3 ;
			RECT 15.761 50.180 16.009 50.260 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[75]

	PIN Q[76]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 50.684 16.009 50.764 ;
			LAYER M2 ;
			RECT 15.761 50.684 16.009 50.764 ;
			LAYER M3 ;
			RECT 15.761 50.684 16.009 50.764 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[76]

	PIN Q[77]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 51.188 16.009 51.268 ;
			LAYER M2 ;
			RECT 15.761 51.188 16.009 51.268 ;
			LAYER M3 ;
			RECT 15.761 51.188 16.009 51.268 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[77]

	PIN Q[78]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 51.692 16.009 51.772 ;
			LAYER M2 ;
			RECT 15.761 51.692 16.009 51.772 ;
			LAYER M3 ;
			RECT 15.761 51.692 16.009 51.772 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[78]

	PIN Q[79]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 52.196 16.009 52.276 ;
			LAYER M2 ;
			RECT 15.761 52.196 16.009 52.276 ;
			LAYER M3 ;
			RECT 15.761 52.196 16.009 52.276 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[79]

	PIN Q[80]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 52.700 16.009 52.780 ;
			LAYER M2 ;
			RECT 15.761 52.700 16.009 52.780 ;
			LAYER M3 ;
			RECT 15.761 52.700 16.009 52.780 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[80]

	PIN Q[81]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 53.204 16.009 53.284 ;
			LAYER M2 ;
			RECT 15.761 53.204 16.009 53.284 ;
			LAYER M3 ;
			RECT 15.761 53.204 16.009 53.284 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[81]

	PIN Q[82]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 53.708 16.009 53.788 ;
			LAYER M2 ;
			RECT 15.761 53.708 16.009 53.788 ;
			LAYER M3 ;
			RECT 15.761 53.708 16.009 53.788 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[82]

	PIN Q[83]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 54.212 16.009 54.292 ;
			LAYER M2 ;
			RECT 15.761 54.212 16.009 54.292 ;
			LAYER M3 ;
			RECT 15.761 54.212 16.009 54.292 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[83]

	PIN Q[84]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 54.716 16.009 54.796 ;
			LAYER M2 ;
			RECT 15.761 54.716 16.009 54.796 ;
			LAYER M3 ;
			RECT 15.761 54.716 16.009 54.796 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[84]

	PIN Q[85]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 55.220 16.009 55.300 ;
			LAYER M2 ;
			RECT 15.761 55.220 16.009 55.300 ;
			LAYER M3 ;
			RECT 15.761 55.220 16.009 55.300 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[85]

	PIN Q[86]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 55.724 16.009 55.804 ;
			LAYER M2 ;
			RECT 15.761 55.724 16.009 55.804 ;
			LAYER M3 ;
			RECT 15.761 55.724 16.009 55.804 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[86]

	PIN Q[87]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 56.228 16.009 56.308 ;
			LAYER M2 ;
			RECT 15.761 56.228 16.009 56.308 ;
			LAYER M3 ;
			RECT 15.761 56.228 16.009 56.308 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[87]

	PIN Q[88]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 56.732 16.009 56.812 ;
			LAYER M2 ;
			RECT 15.761 56.732 16.009 56.812 ;
			LAYER M3 ;
			RECT 15.761 56.732 16.009 56.812 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[88]

	PIN Q[89]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 57.236 16.009 57.316 ;
			LAYER M2 ;
			RECT 15.761 57.236 16.009 57.316 ;
			LAYER M3 ;
			RECT 15.761 57.236 16.009 57.316 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[89]

	PIN Q[90]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 57.740 16.009 57.820 ;
			LAYER M2 ;
			RECT 15.761 57.740 16.009 57.820 ;
			LAYER M3 ;
			RECT 15.761 57.740 16.009 57.820 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[90]

	PIN Q[91]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 58.244 16.009 58.324 ;
			LAYER M2 ;
			RECT 15.761 58.244 16.009 58.324 ;
			LAYER M3 ;
			RECT 15.761 58.244 16.009 58.324 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[91]

	PIN Q[92]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 58.748 16.009 58.828 ;
			LAYER M2 ;
			RECT 15.761 58.748 16.009 58.828 ;
			LAYER M3 ;
			RECT 15.761 58.748 16.009 58.828 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[92]

	PIN Q[93]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 59.252 16.009 59.332 ;
			LAYER M2 ;
			RECT 15.761 59.252 16.009 59.332 ;
			LAYER M3 ;
			RECT 15.761 59.252 16.009 59.332 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[93]

	PIN Q[94]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 59.756 16.009 59.836 ;
			LAYER M2 ;
			RECT 15.761 59.756 16.009 59.836 ;
			LAYER M3 ;
			RECT 15.761 59.756 16.009 59.836 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[94]

	PIN Q[95]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 60.260 16.009 60.340 ;
			LAYER M2 ;
			RECT 15.761 60.260 16.009 60.340 ;
			LAYER M3 ;
			RECT 15.761 60.260 16.009 60.340 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[95]

	PIN Q[96]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 60.764 16.009 60.844 ;
			LAYER M2 ;
			RECT 15.761 60.764 16.009 60.844 ;
			LAYER M3 ;
			RECT 15.761 60.764 16.009 60.844 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[96]

	PIN Q[97]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 61.268 16.009 61.348 ;
			LAYER M2 ;
			RECT 15.761 61.268 16.009 61.348 ;
			LAYER M3 ;
			RECT 15.761 61.268 16.009 61.348 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[97]

	PIN Q[98]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 61.772 16.009 61.852 ;
			LAYER M2 ;
			RECT 15.761 61.772 16.009 61.852 ;
			LAYER M3 ;
			RECT 15.761 61.772 16.009 61.852 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[98]

	PIN Q[99]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 62.276 16.009 62.356 ;
			LAYER M2 ;
			RECT 15.761 62.276 16.009 62.356 ;
			LAYER M3 ;
			RECT 15.761 62.276 16.009 62.356 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[99]

	PIN Q[100]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 62.780 16.009 62.860 ;
			LAYER M2 ;
			RECT 15.761 62.780 16.009 62.860 ;
			LAYER M3 ;
			RECT 15.761 62.780 16.009 62.860 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[100]

	PIN Q[101]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 63.284 16.009 63.364 ;
			LAYER M2 ;
			RECT 15.761 63.284 16.009 63.364 ;
			LAYER M3 ;
			RECT 15.761 63.284 16.009 63.364 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[101]

	PIN Q[102]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 63.788 16.009 63.868 ;
			LAYER M2 ;
			RECT 15.761 63.788 16.009 63.868 ;
			LAYER M3 ;
			RECT 15.761 63.788 16.009 63.868 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[102]

	PIN Q[103]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 64.292 16.009 64.372 ;
			LAYER M2 ;
			RECT 15.761 64.292 16.009 64.372 ;
			LAYER M3 ;
			RECT 15.761 64.292 16.009 64.372 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[103]

	PIN Q[104]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 64.796 16.009 64.876 ;
			LAYER M2 ;
			RECT 15.761 64.796 16.009 64.876 ;
			LAYER M3 ;
			RECT 15.761 64.796 16.009 64.876 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[104]

	PIN Q[105]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 65.300 16.009 65.380 ;
			LAYER M2 ;
			RECT 15.761 65.300 16.009 65.380 ;
			LAYER M3 ;
			RECT 15.761 65.300 16.009 65.380 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[105]

	PIN Q[106]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 65.804 16.009 65.884 ;
			LAYER M2 ;
			RECT 15.761 65.804 16.009 65.884 ;
			LAYER M3 ;
			RECT 15.761 65.804 16.009 65.884 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[106]

	PIN Q[107]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 66.308 16.009 66.388 ;
			LAYER M2 ;
			RECT 15.761 66.308 16.009 66.388 ;
			LAYER M3 ;
			RECT 15.761 66.308 16.009 66.388 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[107]

	PIN Q[108]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 66.812 16.009 66.892 ;
			LAYER M2 ;
			RECT 15.761 66.812 16.009 66.892 ;
			LAYER M3 ;
			RECT 15.761 66.812 16.009 66.892 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[108]

	PIN Q[109]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 67.316 16.009 67.396 ;
			LAYER M2 ;
			RECT 15.761 67.316 16.009 67.396 ;
			LAYER M3 ;
			RECT 15.761 67.316 16.009 67.396 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[109]

	PIN Q[110]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 67.820 16.009 67.900 ;
			LAYER M2 ;
			RECT 15.761 67.820 16.009 67.900 ;
			LAYER M3 ;
			RECT 15.761 67.820 16.009 67.900 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[110]

	PIN Q[111]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 68.324 16.009 68.404 ;
			LAYER M2 ;
			RECT 15.761 68.324 16.009 68.404 ;
			LAYER M3 ;
			RECT 15.761 68.324 16.009 68.404 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[111]

	PIN Q[112]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 68.828 16.009 68.908 ;
			LAYER M2 ;
			RECT 15.761 68.828 16.009 68.908 ;
			LAYER M3 ;
			RECT 15.761 68.828 16.009 68.908 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[112]

	PIN Q[113]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 69.332 16.009 69.412 ;
			LAYER M2 ;
			RECT 15.761 69.332 16.009 69.412 ;
			LAYER M3 ;
			RECT 15.761 69.332 16.009 69.412 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[113]

	PIN Q[114]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 69.836 16.009 69.916 ;
			LAYER M2 ;
			RECT 15.761 69.836 16.009 69.916 ;
			LAYER M3 ;
			RECT 15.761 69.836 16.009 69.916 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[114]

	PIN Q[115]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 70.340 16.009 70.420 ;
			LAYER M2 ;
			RECT 15.761 70.340 16.009 70.420 ;
			LAYER M3 ;
			RECT 15.761 70.340 16.009 70.420 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[115]

	PIN Q[116]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 70.844 16.009 70.924 ;
			LAYER M2 ;
			RECT 15.761 70.844 16.009 70.924 ;
			LAYER M3 ;
			RECT 15.761 70.844 16.009 70.924 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[116]

	PIN Q[117]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 71.348 16.009 71.428 ;
			LAYER M2 ;
			RECT 15.761 71.348 16.009 71.428 ;
			LAYER M3 ;
			RECT 15.761 71.348 16.009 71.428 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[117]

	PIN Q[118]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 71.852 16.009 71.932 ;
			LAYER M2 ;
			RECT 15.761 71.852 16.009 71.932 ;
			LAYER M3 ;
			RECT 15.761 71.852 16.009 71.932 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[118]

	PIN Q[119]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 72.356 16.009 72.436 ;
			LAYER M2 ;
			RECT 15.761 72.356 16.009 72.436 ;
			LAYER M3 ;
			RECT 15.761 72.356 16.009 72.436 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[119]

	PIN Q[120]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 72.860 16.009 72.940 ;
			LAYER M2 ;
			RECT 15.761 72.860 16.009 72.940 ;
			LAYER M3 ;
			RECT 15.761 72.860 16.009 72.940 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[120]

	PIN Q[121]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 73.364 16.009 73.444 ;
			LAYER M2 ;
			RECT 15.761 73.364 16.009 73.444 ;
			LAYER M3 ;
			RECT 15.761 73.364 16.009 73.444 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[121]

	PIN Q[122]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 73.868 16.009 73.948 ;
			LAYER M2 ;
			RECT 15.761 73.868 16.009 73.948 ;
			LAYER M3 ;
			RECT 15.761 73.868 16.009 73.948 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[122]

	PIN Q[123]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 74.372 16.009 74.452 ;
			LAYER M2 ;
			RECT 15.761 74.372 16.009 74.452 ;
			LAYER M3 ;
			RECT 15.761 74.372 16.009 74.452 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[123]

	PIN Q[124]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 74.876 16.009 74.956 ;
			LAYER M2 ;
			RECT 15.761 74.876 16.009 74.956 ;
			LAYER M3 ;
			RECT 15.761 74.876 16.009 74.956 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[124]

	PIN Q[125]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 75.380 16.009 75.460 ;
			LAYER M2 ;
			RECT 15.761 75.380 16.009 75.460 ;
			LAYER M3 ;
			RECT 15.761 75.380 16.009 75.460 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[125]

	PIN Q[126]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 75.884 16.009 75.964 ;
			LAYER M2 ;
			RECT 15.761 75.884 16.009 75.964 ;
			LAYER M3 ;
			RECT 15.761 75.884 16.009 75.964 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[126]

	PIN Q[127]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 76.388 16.009 76.468 ;
			LAYER M2 ;
			RECT 15.761 76.388 16.009 76.468 ;
			LAYER M3 ;
			RECT 15.761 76.388 16.009 76.468 ;
		END
		ANTENNADIFFAREA 0.037083 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.154680 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.009840 LAYER VIA1 ;
		ANTENNADIFFAREA 0.037083 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.163080 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA2 ;
		ANTENNADIFFAREA 0.037083 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.410880 LAYER M3 ;
	END Q[127]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 35.432 16.009 35.512 ;
			LAYER M2 ;
			RECT 15.761 35.432 16.009 35.512 ;
			LAYER M3 ;
			RECT 15.761 35.432 16.009 35.512 ;
		END
		ANTENNAGATEAREA 0.003500 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.087960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.421700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003500 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.054840 LAYER M2 ;
		ANTENNAMAXAREACAR 14.747000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003500 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.753840 LAYER M3 ;
		ANTENNAMAXAREACAR 192.550000 LAYER M3 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 35.816 16.009 35.896 ;
			LAYER M2 ;
			RECT 15.761 35.816 16.009 35.896 ;
			LAYER M3 ;
			RECT 15.761 35.816 16.009 35.896 ;
		END
		ANTENNAGATEAREA 0.003500 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.087960 LAYER M1 ;
		ANTENNAMAXAREACAR 12.421700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003500 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.054840 LAYER M2 ;
		ANTENNAMAXAREACAR 14.747000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003500 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.753840 LAYER M3 ;
		ANTENNAMAXAREACAR 192.550000 LAYER M3 ;
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.176 15.889 1.296 ;
			LAYER M4 ;
			RECT 0.120 1.428 15.889 1.548 ;
			LAYER M4 ;
			RECT 0.120 2.184 15.889 2.304 ;
			LAYER M4 ;
			RECT 0.120 2.436 15.889 2.556 ;
			LAYER M4 ;
			RECT 0.120 3.192 15.889 3.312 ;
			LAYER M4 ;
			RECT 0.120 3.444 15.889 3.564 ;
			LAYER M4 ;
			RECT 0.120 4.200 15.889 4.320 ;
			LAYER M4 ;
			RECT 0.120 4.452 15.889 4.572 ;
			LAYER M4 ;
			RECT 0.120 5.208 15.889 5.328 ;
			LAYER M4 ;
			RECT 0.120 5.460 15.889 5.580 ;
			LAYER M4 ;
			RECT 0.120 6.216 15.889 6.336 ;
			LAYER M4 ;
			RECT 0.120 6.468 15.889 6.588 ;
			LAYER M4 ;
			RECT 0.120 7.224 15.889 7.344 ;
			LAYER M4 ;
			RECT 0.120 7.476 15.889 7.596 ;
			LAYER M4 ;
			RECT 0.120 8.232 15.889 8.352 ;
			LAYER M4 ;
			RECT 0.120 8.484 15.889 8.604 ;
			LAYER M4 ;
			RECT 0.120 9.240 15.889 9.360 ;
			LAYER M4 ;
			RECT 0.120 9.492 15.889 9.612 ;
			LAYER M4 ;
			RECT 0.120 10.248 15.889 10.368 ;
			LAYER M4 ;
			RECT 0.120 10.500 15.889 10.620 ;
			LAYER M4 ;
			RECT 0.120 11.256 15.889 11.376 ;
			LAYER M4 ;
			RECT 0.120 11.508 15.889 11.628 ;
			LAYER M4 ;
			RECT 0.120 12.264 15.889 12.384 ;
			LAYER M4 ;
			RECT 0.120 12.516 15.889 12.636 ;
			LAYER M4 ;
			RECT 0.120 13.272 15.889 13.392 ;
			LAYER M4 ;
			RECT 0.120 13.524 15.889 13.644 ;
			LAYER M4 ;
			RECT 0.120 14.280 15.889 14.400 ;
			LAYER M4 ;
			RECT 0.120 14.532 15.889 14.652 ;
			LAYER M4 ;
			RECT 0.120 15.288 15.889 15.408 ;
			LAYER M4 ;
			RECT 0.120 15.540 15.889 15.660 ;
			LAYER M4 ;
			RECT 0.120 16.296 15.889 16.416 ;
			LAYER M4 ;
			RECT 0.120 16.548 15.889 16.668 ;
			LAYER M4 ;
			RECT 0.120 17.304 15.889 17.424 ;
			LAYER M4 ;
			RECT 0.120 17.556 15.889 17.676 ;
			LAYER M4 ;
			RECT 0.120 18.312 15.889 18.432 ;
			LAYER M4 ;
			RECT 0.120 18.564 15.889 18.684 ;
			LAYER M4 ;
			RECT 0.120 19.320 15.889 19.440 ;
			LAYER M4 ;
			RECT 0.120 19.572 15.889 19.692 ;
			LAYER M4 ;
			RECT 0.120 20.328 15.889 20.448 ;
			LAYER M4 ;
			RECT 0.120 20.580 15.889 20.700 ;
			LAYER M4 ;
			RECT 0.120 21.336 15.889 21.456 ;
			LAYER M4 ;
			RECT 0.120 21.588 15.889 21.708 ;
			LAYER M4 ;
			RECT 0.120 22.344 15.889 22.464 ;
			LAYER M4 ;
			RECT 0.120 22.596 15.889 22.716 ;
			LAYER M4 ;
			RECT 0.120 23.352 15.889 23.472 ;
			LAYER M4 ;
			RECT 0.120 23.604 15.889 23.724 ;
			LAYER M4 ;
			RECT 0.120 24.360 15.889 24.480 ;
			LAYER M4 ;
			RECT 0.120 24.612 15.889 24.732 ;
			LAYER M4 ;
			RECT 0.120 25.368 15.889 25.488 ;
			LAYER M4 ;
			RECT 0.120 25.620 15.889 25.740 ;
			LAYER M4 ;
			RECT 0.120 26.376 15.889 26.496 ;
			LAYER M4 ;
			RECT 0.120 26.628 15.889 26.748 ;
			LAYER M4 ;
			RECT 0.120 27.384 15.889 27.504 ;
			LAYER M4 ;
			RECT 0.120 27.636 15.889 27.756 ;
			LAYER M4 ;
			RECT 0.120 28.392 15.889 28.512 ;
			LAYER M4 ;
			RECT 0.120 28.644 15.889 28.764 ;
			LAYER M4 ;
			RECT 0.120 29.400 15.889 29.520 ;
			LAYER M4 ;
			RECT 0.120 29.652 15.889 29.772 ;
			LAYER M4 ;
			RECT 0.120 30.408 15.889 30.528 ;
			LAYER M4 ;
			RECT 0.120 30.660 15.889 30.780 ;
			LAYER M4 ;
			RECT 0.120 31.416 15.889 31.536 ;
			LAYER M4 ;
			RECT 0.120 31.668 15.889 31.788 ;
			LAYER M4 ;
			RECT 0.120 32.424 15.889 32.544 ;
			LAYER M4 ;
			RECT 0.120 32.676 15.889 32.796 ;
			LAYER M4 ;
			RECT 0.120 34.329 15.889 34.449 ;
			LAYER M4 ;
			RECT 0.120 34.789 15.889 34.909 ;
			LAYER M4 ;
			RECT 0.120 35.249 15.889 35.369 ;
			LAYER M4 ;
			RECT 0.120 35.709 15.889 35.829 ;
			LAYER M4 ;
			RECT 0.120 36.319 15.889 36.439 ;
			LAYER M4 ;
			RECT 0.120 37.009 15.889 37.129 ;
			LAYER M4 ;
			RECT 0.120 37.239 15.889 37.359 ;
			LAYER M4 ;
			RECT 0.120 37.699 15.889 37.819 ;
			LAYER M4 ;
			RECT 0.120 38.159 15.889 38.279 ;
			LAYER M4 ;
			RECT 0.120 38.739 15.889 38.859 ;
			LAYER M4 ;
			RECT 0.120 39.429 15.889 39.549 ;
			LAYER M4 ;
			RECT 0.120 39.659 15.889 39.779 ;
			LAYER M4 ;
			RECT 0.120 39.889 15.889 40.009 ;
			LAYER M4 ;
			RECT 0.120 40.964 15.889 41.084 ;
			LAYER M4 ;
			RECT 0.120 41.819 15.889 41.939 ;
			LAYER M4 ;
			RECT 0.120 42.279 15.889 42.399 ;
			LAYER M4 ;
			RECT 0.120 42.739 15.889 42.859 ;
			LAYER M4 ;
			RECT 0.120 43.589 15.889 43.709 ;
			LAYER M4 ;
			RECT 0.120 44.616 15.889 44.736 ;
			LAYER M4 ;
			RECT 0.120 44.868 15.889 44.988 ;
			LAYER M4 ;
			RECT 0.120 45.624 15.889 45.744 ;
			LAYER M4 ;
			RECT 0.120 45.876 15.889 45.996 ;
			LAYER M4 ;
			RECT 0.120 46.632 15.889 46.752 ;
			LAYER M4 ;
			RECT 0.120 46.884 15.889 47.004 ;
			LAYER M4 ;
			RECT 0.120 47.640 15.889 47.760 ;
			LAYER M4 ;
			RECT 0.120 47.892 15.889 48.012 ;
			LAYER M4 ;
			RECT 0.120 48.648 15.889 48.768 ;
			LAYER M4 ;
			RECT 0.120 48.900 15.889 49.020 ;
			LAYER M4 ;
			RECT 0.120 49.656 15.889 49.776 ;
			LAYER M4 ;
			RECT 0.120 49.908 15.889 50.028 ;
			LAYER M4 ;
			RECT 0.120 50.664 15.889 50.784 ;
			LAYER M4 ;
			RECT 0.120 50.916 15.889 51.036 ;
			LAYER M4 ;
			RECT 0.120 51.672 15.889 51.792 ;
			LAYER M4 ;
			RECT 0.120 51.924 15.889 52.044 ;
			LAYER M4 ;
			RECT 0.120 52.680 15.889 52.800 ;
			LAYER M4 ;
			RECT 0.120 52.932 15.889 53.052 ;
			LAYER M4 ;
			RECT 0.120 53.688 15.889 53.808 ;
			LAYER M4 ;
			RECT 0.120 53.940 15.889 54.060 ;
			LAYER M4 ;
			RECT 0.120 54.696 15.889 54.816 ;
			LAYER M4 ;
			RECT 0.120 54.948 15.889 55.068 ;
			LAYER M4 ;
			RECT 0.120 55.704 15.889 55.824 ;
			LAYER M4 ;
			RECT 0.120 55.956 15.889 56.076 ;
			LAYER M4 ;
			RECT 0.120 56.712 15.889 56.832 ;
			LAYER M4 ;
			RECT 0.120 56.964 15.889 57.084 ;
			LAYER M4 ;
			RECT 0.120 57.720 15.889 57.840 ;
			LAYER M4 ;
			RECT 0.120 57.972 15.889 58.092 ;
			LAYER M4 ;
			RECT 0.120 58.728 15.889 58.848 ;
			LAYER M4 ;
			RECT 0.120 58.980 15.889 59.100 ;
			LAYER M4 ;
			RECT 0.120 59.736 15.889 59.856 ;
			LAYER M4 ;
			RECT 0.120 59.988 15.889 60.108 ;
			LAYER M4 ;
			RECT 0.120 60.744 15.889 60.864 ;
			LAYER M4 ;
			RECT 0.120 60.996 15.889 61.116 ;
			LAYER M4 ;
			RECT 0.120 61.752 15.889 61.872 ;
			LAYER M4 ;
			RECT 0.120 62.004 15.889 62.124 ;
			LAYER M4 ;
			RECT 0.120 62.760 15.889 62.880 ;
			LAYER M4 ;
			RECT 0.120 63.012 15.889 63.132 ;
			LAYER M4 ;
			RECT 0.120 63.768 15.889 63.888 ;
			LAYER M4 ;
			RECT 0.120 64.020 15.889 64.140 ;
			LAYER M4 ;
			RECT 0.120 64.776 15.889 64.896 ;
			LAYER M4 ;
			RECT 0.120 65.028 15.889 65.148 ;
			LAYER M4 ;
			RECT 0.120 65.784 15.889 65.904 ;
			LAYER M4 ;
			RECT 0.120 66.036 15.889 66.156 ;
			LAYER M4 ;
			RECT 0.120 66.792 15.889 66.912 ;
			LAYER M4 ;
			RECT 0.120 67.044 15.889 67.164 ;
			LAYER M4 ;
			RECT 0.120 67.800 15.889 67.920 ;
			LAYER M4 ;
			RECT 0.120 68.052 15.889 68.172 ;
			LAYER M4 ;
			RECT 0.120 68.808 15.889 68.928 ;
			LAYER M4 ;
			RECT 0.120 69.060 15.889 69.180 ;
			LAYER M4 ;
			RECT 0.120 69.816 15.889 69.936 ;
			LAYER M4 ;
			RECT 0.120 70.068 15.889 70.188 ;
			LAYER M4 ;
			RECT 0.120 70.824 15.889 70.944 ;
			LAYER M4 ;
			RECT 0.120 71.076 15.889 71.196 ;
			LAYER M4 ;
			RECT 0.120 71.832 15.889 71.952 ;
			LAYER M4 ;
			RECT 0.120 72.084 15.889 72.204 ;
			LAYER M4 ;
			RECT 0.120 72.840 15.889 72.960 ;
			LAYER M4 ;
			RECT 0.120 73.092 15.889 73.212 ;
			LAYER M4 ;
			RECT 0.120 73.848 15.889 73.968 ;
			LAYER M4 ;
			RECT 0.120 74.100 15.889 74.220 ;
			LAYER M4 ;
			RECT 0.120 74.856 15.889 74.976 ;
			LAYER M4 ;
			RECT 0.120 75.108 15.889 75.228 ;
			LAYER M4 ;
			RECT 0.120 75.864 15.889 75.984 ;
			LAYER M4 ;
			RECT 0.120 76.116 15.889 76.236 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 0.321 15.889 0.481 ;
			LAYER M4 ;
			RECT 0.120 0.924 15.889 1.044 ;
			LAYER M4 ;
			RECT 0.120 1.932 15.889 2.052 ;
			LAYER M4 ;
			RECT 0.120 2.940 15.889 3.060 ;
			LAYER M4 ;
			RECT 0.120 3.948 15.889 4.068 ;
			LAYER M4 ;
			RECT 0.120 4.956 15.889 5.076 ;
			LAYER M4 ;
			RECT 0.120 5.964 15.889 6.084 ;
			LAYER M4 ;
			RECT 0.120 6.972 15.889 7.092 ;
			LAYER M4 ;
			RECT 0.120 7.980 15.889 8.100 ;
			LAYER M4 ;
			RECT 0.120 8.988 15.889 9.108 ;
			LAYER M4 ;
			RECT 0.120 9.996 15.889 10.116 ;
			LAYER M4 ;
			RECT 0.120 11.004 15.889 11.124 ;
			LAYER M4 ;
			RECT 0.120 12.012 15.889 12.132 ;
			LAYER M4 ;
			RECT 0.120 13.020 15.889 13.140 ;
			LAYER M4 ;
			RECT 0.120 14.028 15.889 14.148 ;
			LAYER M4 ;
			RECT 0.120 15.036 15.889 15.156 ;
			LAYER M4 ;
			RECT 0.120 16.044 15.889 16.164 ;
			LAYER M4 ;
			RECT 0.120 17.052 15.889 17.172 ;
			LAYER M4 ;
			RECT 0.120 18.060 15.889 18.180 ;
			LAYER M4 ;
			RECT 0.120 19.068 15.889 19.188 ;
			LAYER M4 ;
			RECT 0.120 20.076 15.889 20.196 ;
			LAYER M4 ;
			RECT 0.120 21.084 15.889 21.204 ;
			LAYER M4 ;
			RECT 0.120 22.092 15.889 22.212 ;
			LAYER M4 ;
			RECT 0.120 23.100 15.889 23.220 ;
			LAYER M4 ;
			RECT 0.120 24.108 15.889 24.228 ;
			LAYER M4 ;
			RECT 0.120 25.116 15.889 25.236 ;
			LAYER M4 ;
			RECT 0.120 26.124 15.889 26.244 ;
			LAYER M4 ;
			RECT 0.120 27.132 15.889 27.252 ;
			LAYER M4 ;
			RECT 0.120 28.140 15.889 28.260 ;
			LAYER M4 ;
			RECT 0.120 29.148 15.889 29.268 ;
			LAYER M4 ;
			RECT 0.120 30.156 15.889 30.276 ;
			LAYER M4 ;
			RECT 0.120 31.164 15.889 31.284 ;
			LAYER M4 ;
			RECT 0.120 32.172 15.889 32.292 ;
			LAYER M4 ;
			RECT 0.120 33.180 15.889 33.300 ;
			LAYER M4 ;
			RECT 0.120 34.559 15.889 34.679 ;
			LAYER M4 ;
			RECT 0.120 35.019 15.889 35.139 ;
			LAYER M4 ;
			RECT 0.120 35.479 15.889 35.599 ;
			LAYER M4 ;
			RECT 0.120 36.089 15.889 36.209 ;
			LAYER M4 ;
			RECT 0.120 36.549 15.889 36.669 ;
			LAYER M4 ;
			RECT 0.120 36.779 15.889 36.899 ;
			LAYER M4 ;
			RECT 0.120 37.469 15.889 37.589 ;
			LAYER M4 ;
			RECT 0.120 37.929 15.889 38.049 ;
			LAYER M4 ;
			RECT 0.120 38.509 15.889 38.629 ;
			LAYER M4 ;
			RECT 0.120 38.969 15.889 39.089 ;
			LAYER M4 ;
			RECT 0.120 39.199 15.889 39.319 ;
			LAYER M4 ;
			RECT 0.120 40.119 15.889 40.239 ;
			LAYER M4 ;
			RECT 0.120 40.504 15.889 40.624 ;
			LAYER M4 ;
			RECT 0.120 40.734 15.889 40.854 ;
			LAYER M4 ;
			RECT 0.120 41.194 15.889 41.314 ;
			LAYER M4 ;
			RECT 0.120 41.589 15.889 41.709 ;
			LAYER M4 ;
			RECT 0.120 42.049 15.889 42.169 ;
			LAYER M4 ;
			RECT 0.120 42.509 15.889 42.629 ;
			LAYER M4 ;
			RECT 0.120 42.969 15.889 43.089 ;
			LAYER M4 ;
			RECT 0.120 43.359 15.889 43.479 ;
			LAYER M4 ;
			RECT 0.120 43.819 15.889 43.939 ;
			LAYER M4 ;
			RECT 0.120 44.364 15.889 44.484 ;
			LAYER M4 ;
			RECT 0.120 45.372 15.889 45.492 ;
			LAYER M4 ;
			RECT 0.120 46.380 15.889 46.500 ;
			LAYER M4 ;
			RECT 0.120 47.388 15.889 47.508 ;
			LAYER M4 ;
			RECT 0.120 48.396 15.889 48.516 ;
			LAYER M4 ;
			RECT 0.120 49.404 15.889 49.524 ;
			LAYER M4 ;
			RECT 0.120 50.412 15.889 50.532 ;
			LAYER M4 ;
			RECT 0.120 51.420 15.889 51.540 ;
			LAYER M4 ;
			RECT 0.120 52.428 15.889 52.548 ;
			LAYER M4 ;
			RECT 0.120 53.436 15.889 53.556 ;
			LAYER M4 ;
			RECT 0.120 54.444 15.889 54.564 ;
			LAYER M4 ;
			RECT 0.120 55.452 15.889 55.572 ;
			LAYER M4 ;
			RECT 0.120 56.460 15.889 56.580 ;
			LAYER M4 ;
			RECT 0.120 57.468 15.889 57.588 ;
			LAYER M4 ;
			RECT 0.120 58.476 15.889 58.596 ;
			LAYER M4 ;
			RECT 0.120 59.484 15.889 59.604 ;
			LAYER M4 ;
			RECT 0.120 60.492 15.889 60.612 ;
			LAYER M4 ;
			RECT 0.120 61.500 15.889 61.620 ;
			LAYER M4 ;
			RECT 0.120 62.508 15.889 62.628 ;
			LAYER M4 ;
			RECT 0.120 63.516 15.889 63.636 ;
			LAYER M4 ;
			RECT 0.120 64.524 15.889 64.644 ;
			LAYER M4 ;
			RECT 0.120 65.532 15.889 65.652 ;
			LAYER M4 ;
			RECT 0.120 66.540 15.889 66.660 ;
			LAYER M4 ;
			RECT 0.120 67.548 15.889 67.668 ;
			LAYER M4 ;
			RECT 0.120 68.556 15.889 68.676 ;
			LAYER M4 ;
			RECT 0.120 69.564 15.889 69.684 ;
			LAYER M4 ;
			RECT 0.120 70.572 15.889 70.692 ;
			LAYER M4 ;
			RECT 0.120 71.580 15.889 71.700 ;
			LAYER M4 ;
			RECT 0.120 72.588 15.889 72.708 ;
			LAYER M4 ;
			RECT 0.120 73.596 15.889 73.716 ;
			LAYER M4 ;
			RECT 0.120 74.604 15.889 74.724 ;
			LAYER M4 ;
			RECT 0.120 75.612 15.889 75.732 ;
			LAYER M4 ;
			RECT 0.120 76.620 15.889 76.740 ;
			LAYER M4 ;
			RECT 0.120 77.183 15.889 77.343 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 39.464 16.009 39.544 ;
			LAYER M2 ;
			RECT 15.761 39.464 16.009 39.544 ;
			LAYER M3 ;
			RECT 15.761 39.464 16.009 39.544 ;
		END
		ANTENNAGATEAREA 0.001917 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.049680 LAYER M1 ;
		ANTENNAMAXAREACAR 3.793440 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.001917 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.111480 LAYER M2 ;
		ANTENNAMAXAREACAR 16.918900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.001917 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.699360 LAYER M3 ;
		ANTENNAMAXAREACAR 82.231100 LAYER M3 ;
	END WEB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 34.664 16.009 34.744 ;
			LAYER M2 ;
			RECT 15.761 34.664 16.009 34.744 ;
			LAYER M3 ;
			RECT 15.761 34.664 16.009 34.744 ;
		END
		ANTENNAGATEAREA 0.003500 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.104280 LAYER M1 ;
		ANTENNAMAXAREACAR 16.293400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003500 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.073320 LAYER M2 ;
		ANTENNAMAXAREACAR 25.874200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003500 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.746400 LAYER M3 ;
		ANTENNAMAXAREACAR 201.916000 LAYER M3 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.761 35.624 16.009 35.704 ;
			LAYER M2 ;
			RECT 15.761 35.624 16.009 35.704 ;
			LAYER M3 ;
			RECT 15.761 35.624 16.009 35.704 ;
		END
		ANTENNAGATEAREA 0.003500 LAYER M1 ;
		ANTENNADIFFAREA 0.006750 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.104280 LAYER M1 ;
		ANTENNAMAXAREACAR 16.293400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.289800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.003500 LAYER M2 ;
		ANTENNADIFFAREA 0.006750 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.073320 LAYER M2 ;
		ANTENNAMAXAREACAR 25.874200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.579600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.003500 LAYER M3 ;
		ANTENNADIFFAREA 0.006750 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.746400 LAYER M3 ;
		ANTENNAMAXAREACAR 201.916000 LAYER M3 ;
	END WTSEL[1]

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 16.009 77.664 ;
		LAYER M2 ;
		RECT 0.000 0.000 16.009 77.664 ;
		LAYER M3 ;
		RECT 0.000 0.000 16.009 77.664 ;
		LAYER M4 ;
		RECT 0.761 38.290 4.123 38.354 ;
		LAYER M4 ;
		RECT 0.761 40.412 4.303 40.476 ;
		LAYER M4 ;
		RECT 0.761 41.406 4.573 41.470 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 16.009 77.664 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 16.009 77.664 ;
	END
END TS5N16FFCLLSVTA8X128M1SW

END LIBRARY
