**** Created by MC2: Version 2013.12.00.f on 2025/06/23, 09:41:45 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  n16ff_uhd1prf_sb_leafcell
* Top Cell Name: COMPILER_LEAFCELL
* View Name:     schematic
* Netlisted on:  Sep 11 17:24:04 2015
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM


*.PIN vss

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_inv_lvt_mac_pcell_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_lvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_nor2_lvt_mac_pcell_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_lvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_nand3_lvt_mac_pcell_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    MCB_D0907
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_MCB_D0907 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
MNCHPG1 TSMC_2 TSMC_6 TSMC_7 TSMC_5 nchpg_hcsr_mac l=20n nfin=2 m=1 
MNCHPG0 TSMC_1 TSMC_6 TSMC_8 TSMC_5 nchpg_hcsr_mac l=20n nfin=2 m=1 
MNCHPD1 TSMC_7 TSMC_8 TSMC_5 TSMC_5 nchpd_hcsr_mac l=20n nfin=2 m=1 
MNCHPD0 TSMC_8 TSMC_7 TSMC_5 TSMC_5 nchpd_hcsr_mac l=20n nfin=2 m=1 
MPCHPU1 TSMC_7 TSMC_8 TSMC_3 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
MPCHPU0 TSMC_8 TSMC_7 TSMC_3 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    MCB_D0907_ONCELL
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_MCB_D0907_ONCELL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
Mpg11 TSMC_1 TSMC_2 TSMC_9 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd11 TSMC_9 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg21 TSMC_11 TSMC_7 TSMC_10 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_12 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_13 TSMC_12 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_12 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_11 TSMC_8 TSMC_13 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpu11 TSMC_9 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_12 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    WLDRV4X1_core
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_WLDRV4X1_core TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
MM100 TSMC_13 TSMC_17 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM43 TSMC_12 TSMC_18 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM91 TSMC_11 TSMC_19 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM97 TSMC_14 TSMC_20 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM92 TSMC_15 TSMC_19 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM99 TSMC_9 TSMC_17 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM89 TSMC_16 TSMC_18 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM98 TSMC_10 TSMC_20 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=14 m=2 
MM100_2 TSMC_13 TSMC_17 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM43_2 TSMC_12 TSMC_18 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM91_2 TSMC_11 TSMC_19 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM97_2 TSMC_14 TSMC_20 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM92_2 TSMC_15 TSMC_19 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM99_2 TSMC_9 TSMC_17 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM89_2 TSMC_16 TSMC_18 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM98_2 TSMC_10 TSMC_20 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=4 m=2 
MM42 TSMC_12 TSMC_18 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM93 TSMC_11 TSMC_19 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM113 TSMC_21 TSMC_8 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=3 m=4 
MM95 TSMC_14 TSMC_20 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM88 TSMC_22 TSMC_21 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=6 m=8 
MM112 TSMC_21 TSMC_7 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=3 m=4 
MM94 TSMC_15 TSMC_19 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM96 TSMC_10 TSMC_20 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM90 TSMC_16 TSMC_18 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM101 TSMC_9 TSMC_17 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM102 TSMC_13 TSMC_17 TSMC_2 TSMC_2 nch_svt_mac l=20n nfin=12 m=2 
MM79 TSMC_19 TSMC_5 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM82 TSMC_20 TSMC_4 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM85 TSMC_17 TSMC_3 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM18 TSMC_18 TSMC_6 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM111 TSMC_21 TSMC_7 TSMC_23 TSMC_1 pch_lvt_mac l=20n nfin=5 m=4 
MM110 TSMC_23 TSMC_8 TSMC_1 TSMC_1 pch_lvt_mac l=20n nfin=5 m=4 
MM80 TSMC_19 TSMC_21 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM86 TSMC_17 TSMC_21 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM76 TSMC_22 TSMC_21 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=2 m=4 
MM77 TSMC_18 TSMC_21 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM81 TSMC_20 TSMC_21 TSMC_1 TSMC_1 pch_svt_mac l=16.0n nfin=6 m=1 
MM87 TSMC_20 TSMC_4 TSMC_22 TSMC_2 nch_lvt_mac l=16.0n nfin=12 m=1 
MM78 TSMC_19 TSMC_5 TSMC_22 TSMC_2 nch_lvt_mac l=16.0n nfin=12 m=1 
MM84 TSMC_17 TSMC_3 TSMC_22 TSMC_2 nch_lvt_mac l=16.0n nfin=12 m=1 
MM17 TSMC_18 TSMC_6 TSMC_22 TSMC_2 nch_lvt_mac l=16.0n nfin=12 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    WLDRV4X1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_WLDRV4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
XWLDV TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ S5LLSVTSW8U80_WLDRV4X1_core 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_lvt_mac_pcell_4
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    DINB1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_DINB1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 
MM35 TSMC_12 TSMC_13 TSMC_14 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
MM32 TSMC_5 TSMC_7 TSMC_15 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
MM30 TSMC_15 TSMC_16 TSMC_14 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
MM34 TSMC_4 TSMC_7 TSMC_12 TSMC_11 nch_lvt_mac l=20n nfin=3 m=1 
MM33 TSMC_14 TSMC_17 TSMC_11 TSMC_11 nch_lvt_mac l=20n nfin=3 m=2 
MM2 TSMC_18 TSMC_19 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=2 m=2 
MM0 TSMC_16 TSMC_3 TSMC_18 TSMC_11 nch_svt_mac l=20n nfin=2 m=2 
MTN3 TSMC_17 TSMC_1 TSMC_20 TSMC_11 nch_svt_mac l=20n nfin=2 m=2 
MM13 TSMC_17 TSMC_21 TSMC_22 TSMC_11 nch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_23 TSMC_13 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_16 TSMC_21 TSMC_23 TSMC_11 nch_svt_mac l=20n nfin=2 m=1 
MM11 TSMC_22 TSMC_24 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=2 m=1 
MTN2 TSMC_20 TSMC_19 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=2 m=2 
MM29 TSMC_5 TSMC_7 TSMC_10 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MM31 TSMC_5 TSMC_16 TSMC_10 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MM36 TSMC_5 TSMC_17 TSMC_10 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MM37 TSMC_4 TSMC_17 TSMC_10 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MM38 TSMC_4 TSMC_13 TSMC_10 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MM39 TSMC_4 TSMC_7 TSMC_10 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_25 TSMC_21 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=2 m=2 
MM6 TSMC_16 TSMC_3 TSMC_25 TSMC_8 pch_svt_mac l=20n nfin=2 m=2 
MP0 TSMC_26 TSMC_21 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=2 m=2 
MP3 TSMC_17 TSMC_19 TSMC_27 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MP2 TSMC_27 TSMC_24 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MP1 TSMC_17 TSMC_1 TSMC_26 TSMC_8 pch_svt_mac l=20n nfin=2 m=2 
MM3 TSMC_28 TSMC_13 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_16 TSMC_19 TSMC_28 TSMC_8 pch_svt_mac l=20n nfin=2 m=1 
XI66 TSMC_11 TSMC_11 TSMC_24 TSMC_2 TSMC_9 TSMC_8 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI52 TSMC_11 TSMC_11 TSMC_17 TSMC_24 TSMC_9 TSMC_8 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI38 TSMC_11 TSMC_11 TSMC_6 TSMC_19 TSMC_9 TSMC_8 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI18 TSMC_11 TSMC_11 TSMC_16 TSMC_13 TSMC_9 TSMC_8 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI64 TSMC_11 TSMC_11 TSMC_19 TSMC_21 TSMC_9 TSMC_8 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    IOEDGE_R
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_IOEDGE_R TSMC_1 TSMC_2 TSMC_3 TSMC_4 
MM52 TSMC_4 TSMC_1 TSMC_4 TSMC_4 nch_svt_mac l=20n nfin=2 m=1 
MM51 TSMC_2 TSMC_1 TSMC_2 TSMC_2 pch_svt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    DIOB1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_DIOB1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
MM5 TSMC_8 TSMC_7 TSMC_12 TSMC_10 pch_lvt_mac l=20n nfin=3 m=2 
MMP50 TSMC_7 TSMC_9 TSMC_12 TSMC_10 pch_lvt_mac l=20n nfin=3 m=2 
MP1 TSMC_14 TSMC_1 TSMC_11 TSMC_10 pch_ulvt_mac l=20n nfin=4 m=2 
MM0 TSMC_5 TSMC_8 TSMC_14 TSMC_10 pch_ulvt_mac l=20n nfin=4 m=2 
MM3 TSMC_15 TSMC_2 TSMC_11 TSMC_10 pch_ulvt_mac l=20n nfin=4 m=2 
MM4 TSMC_6 TSMC_8 TSMC_15 TSMC_10 pch_ulvt_mac l=20n nfin=4 m=2 
MN1 TSMC_16 TSMC_1 TSMC_13 TSMC_13 nch_svt_mac l=20n nfin=3 m=2 
MM9 TSMC_5 TSMC_7 TSMC_16 TSMC_13 nch_svt_mac l=20n nfin=3 m=2 
MM1 TSMC_6 TSMC_7 TSMC_17 TSMC_13 nch_svt_mac l=20n nfin=3 m=2 
MMN50 TSMC_7 TSMC_9 TSMC_13 TSMC_13 nch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_17 TSMC_2 TSMC_13 TSMC_13 nch_svt_mac l=20n nfin=3 m=2 
MM8 TSMC_8 TSMC_7 TSMC_13 TSMC_13 nch_svt_mac l=20n nfin=3 m=2 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    DOUT1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_DOUT1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
MM6 TSMC_2 TSMC_1 TSMC_6 TSMC_5 pch_svt_mac l=20n nfin=3 m=5 
MM2 TSMC_8 TSMC_9 TSMC_6 TSMC_5 pch_svt_mac l=20n nfin=2 m=1 
MM0 TSMC_1 TSMC_3 TSMC_8 TSMC_5 pch_svt_mac l=20n nfin=2 m=1 
XI30 TSMC_7 TSMC_7 TSMC_1 TSMC_9 TSMC_6 TSMC_5 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
MM7 TSMC_2 TSMC_1 TSMC_7 TSMC_7 nch_svt_mac l=20n nfin=3 m=5 
MM1 TSMC_1 TSMC_4 TSMC_10 TSMC_7 nch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_10 TSMC_9 TSMC_7 TSMC_7 nch_svt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    WRITE_PASS1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_WRITE_PASS1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 
MM21 TSMC_8 TSMC_4 TSMC_7 TSMC_7 nch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_9 TSMC_3 TSMC_7 TSMC_7 nch_svt_mac l=20n nfin=2 m=1 
MN2 TSMC_1 TSMC_8 TSMC_7 TSMC_7 nch_svt_mac l=16n nfin=4 m=2 
MN3 TSMC_2 TSMC_9 TSMC_7 TSMC_7 nch_svt_mac l=16n nfin=4 m=2 
MM10 TSMC_9 TSMC_3 TSMC_6 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MM23 TSMC_8 TSMC_4 TSMC_6 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MM0 TSMC_2 TSMC_4 TSMC_6 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
MM14 TSMC_1 TSMC_3 TSMC_6 TSMC_5 pch_lvt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    SA_MUX1_L20X2
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_SA_MUX1_L20X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 
MM10 TSMC_4 TSMC_11 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=4 m=2 
MM12 TSMC_4 TSMC_2 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=4 m=1 
MM14 TSMC_9 TSMC_11 TSMC_2 TSMC_8 pch_svt_mac l=20n nfin=4 m=2 
MP7 TSMC_9 TSMC_3 TSMC_1 TSMC_8 pch_svt_mac l=20n nfin=4 m=1 
MP2_MIXV_SSS TSMC_9 TSMC_11 TSMC_1 TSMC_8 pch_svt_mac l=20n nfin=4 m=2 
MP6 TSMC_3 TSMC_1 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=4 m=1 
MM8 TSMC_3 TSMC_11 TSMC_1 TSMC_8 pch_svt_mac l=20n nfin=4 m=1 
MM13 TSMC_4 TSMC_11 TSMC_2 TSMC_8 pch_svt_mac l=20n nfin=4 m=1 
MM15 TSMC_9 TSMC_4 TSMC_2 TSMC_8 pch_svt_mac l=20n nfin=4 m=1 
MP3_MIXV_SSS TSMC_3 TSMC_11 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=4 m=2 
XI81 TSMC_6 TSMC_7 TSMC_10 TSMC_10 TSMC_9 TSMC_8 TSMC_11 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=7 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
MM4_MIXV_SSS TSMC_3 TSMC_1 TSMC_12 TSMC_10 nch_svt_mac l=20n nfin=5 m=4 
MM16 TSMC_2 TSMC_4 TSMC_13 TSMC_10 nch_svt_mac l=20n nfin=5 m=4 
MM11 TSMC_4 TSMC_2 TSMC_13 TSMC_10 nch_svt_mac l=20n nfin=5 m=4 
MM2 TSMC_12 TSMC_5 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=5 m=4 
MM17 TSMC_13 TSMC_5 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=5 m=4 
MM10_MIXV_SSS TSMC_1 TSMC_3 TSMC_12 TSMC_10 nch_svt_mac l=20n nfin=5 
+ m=4 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    BIT1A_CORE_L20
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_BIT1A_CORE_L20 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 
Xdiob TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_15 
+ TSMC_18 TSMC_19 TSMC_19 TSMC_21 S5LLSVTSW8U80_DIOB1 
Xdout<0> TSMC_22 TSMC_13 TSMC_24 TSMC_25 TSMC_18 TSMC_19 TSMC_21 
+ S5LLSVTSW8U80_DOUT1 
Xdout<1> TSMC_23 TSMC_14 TSMC_24 TSMC_25 TSMC_18 TSMC_19 TSMC_21 
+ S5LLSVTSW8U80_DOUT1 
Xdinb<0> TSMC_5 TSMC_7 TSMC_9 TSMC_26 TSMC_27 TSMC_11 TSMC_12 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 S5LLSVTSW8U80_DINB1 
Xdinb<1> TSMC_6 TSMC_8 TSMC_10 TSMC_28 TSMC_29 TSMC_11 TSMC_12 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 S5LLSVTSW8U80_DINB1 
Xwpass<0> TSMC_1 TSMC_3 TSMC_26 TSMC_27 TSMC_18 TSMC_20 TSMC_21 
+ S5LLSVTSW8U80_WRITE_PASS1 
Xwpass<1> TSMC_2 TSMC_4 TSMC_28 TSMC_29 TSMC_18 TSMC_20 TSMC_21 
+ S5LLSVTSW8U80_WRITE_PASS1 
XSA<0> TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_24 TSMC_25 TSMC_17 TSMC_18 TSMC_20 
+ TSMC_21 S5LLSVTSW8U80_SA_MUX1_L20X2 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    RESETD_RTSEL
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_RESETD_RTSEL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM24 TSMC_9 TSMC_8 TSMC_6 TSMC_6 nch_svt_mac l=16.0n nfin=2 m=1 
MM8 TSMC_10 TSMC_11 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=2 m=1 
MM19 TSMC_2 TSMC_12 TSMC_9 TSMC_6 nch_svt_mac l=16.0n nfin=2 m=1 
MM6 TSMC_13 TSMC_11 TSMC_10 TSMC_6 nch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_14 TSMC_1 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=2 m=1 
MM2 TSMC_11 TSMC_1 TSMC_14 TSMC_6 nch_svt_mac l=20n nfin=2 m=1 
MM10 TSMC_15 TSMC_13 TSMC_16 TSMC_6 nch_svt_mac l=20n nfin=2 m=1 
MM12 TSMC_16 TSMC_13 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_12 TSMC_17 TSMC_5 TSMC_4 pch_svt_mac l=16.0n nfin=2 m=1 
MM17 TSMC_12 TSMC_1 TSMC_5 TSMC_4 pch_svt_mac l=16.0n nfin=2 m=1 
MM7 TSMC_13 TSMC_11 TSMC_18 TSMC_4 pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_19 TSMC_1 TSMC_5 TSMC_4 pch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_11 TSMC_1 TSMC_19 TSMC_4 pch_svt_mac l=20n nfin=2 m=1 
MM9 TSMC_18 TSMC_11 TSMC_5 TSMC_4 pch_svt_mac l=20n nfin=2 m=1 
MM11 TSMC_15 TSMC_13 TSMC_20 TSMC_4 pch_svt_mac l=20n nfin=2 m=1 
MM13 TSMC_20 TSMC_13 TSMC_5 TSMC_4 pch_svt_mac l=20n nfin=2 m=1 
XI8 TSMC_6 TSMC_6 TSMC_7 TSMC_21 TSMC_5 TSMC_4 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI7 TSMC_6 TSMC_6 TSMC_8 TSMC_22 TSMC_5 TSMC_4 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI14 TSMC_7 TSMC_8 TSMC_6 TSMC_6 TSMC_5 TSMC_4 TSMC_23 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI0 TSMC_23 TSMC_15 TSMC_6 TSMC_6 TSMC_5 TSMC_4 TSMC_24 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI11 TSMC_1 TSMC_24 TSMC_6 TSMC_6 TSMC_5 TSMC_4 TSMC_25 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI10 TSMC_25 TSMC_26 TSMC_6 TSMC_6 TSMC_5 TSMC_4 TSMC_17 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI12 TSMC_21 TSMC_8 TSMC_6 TSMC_6 TSMC_5 TSMC_4 TSMC_26 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
MM14 TSMC_27 TSMC_17 TSMC_6 TSMC_6 nch_ulvt_mac l=16.0n nfin=2 m=1 
MM15 TSMC_12 TSMC_1 TSMC_27 TSMC_6 nch_ulvt_mac l=16.0n nfin=2 m=1 
MM23 TSMC_2 TSMC_8 TSMC_5 TSMC_4 pch_ulvt_mac l=16.0n nfin=6 m=1 
MM21 TSMC_2 TSMC_12 TSMC_5 TSMC_4 pch_ulvt_mac l=16.0n nfin=6 m=1 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_ulvt_mac_pcell_6
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_nand3_ulvt_mac_pcell_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    RESETD_WTSEL
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_RESETD_WTSEL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM8 TSMC_9 TSMC_10 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=2 m=1 
MM6 TSMC_11 TSMC_10 TSMC_9 TSMC_5 nch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_12 TSMC_1 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=2 m=1 
MM2 TSMC_10 TSMC_1 TSMC_12 TSMC_5 nch_svt_mac l=20n nfin=2 m=1 
MM10 TSMC_13 TSMC_11 TSMC_14 TSMC_5 nch_svt_mac l=20n nfin=2 m=1 
MM12 TSMC_14 TSMC_11 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=2 m=1 
MM20 TSMC_15 TSMC_1 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM18 TSMC_16 TSMC_17 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM17 TSMC_16 TSMC_18 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_11 TSMC_10 TSMC_19 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM19 TSMC_15 TSMC_20 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_21 TSMC_1 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_10 TSMC_1 TSMC_21 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM9 TSMC_19 TSMC_10 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM11 TSMC_13 TSMC_11 TSMC_22 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
MM13 TSMC_22 TSMC_11 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=2 m=1 
XI8 TSMC_5 TSMC_5 TSMC_7 TSMC_17 TSMC_4 TSMC_3 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI7 TSMC_5 TSMC_5 TSMC_8 TSMC_18 TSMC_4 TSMC_3 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI14 TSMC_17 TSMC_8 TSMC_5 TSMC_5 TSMC_4 TSMC_3 TSMC_23 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI0 TSMC_23 TSMC_13 TSMC_5 TSMC_5 TSMC_4 TSMC_3 TSMC_24 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI11 TSMC_1 TSMC_24 TSMC_5 TSMC_5 TSMC_4 TSMC_3 TSMC_25 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI10 TSMC_25 TSMC_26 TSMC_5 TSMC_5 TSMC_4 TSMC_3 TSMC_20 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI12 TSMC_7 TSMC_18 TSMC_5 TSMC_5 TSMC_4 TSMC_3 TSMC_26 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
MM0 TSMC_16 TSMC_17 TSMC_27 TSMC_5 nch_ulvt_mac l=20n nfin=2 m=1 
MM1 TSMC_27 TSMC_18 TSMC_5 TSMC_5 nch_ulvt_mac l=20n nfin=2 m=1 
MM15 TSMC_15 TSMC_1 TSMC_28 TSMC_5 nch_ulvt_mac l=20n nfin=2 m=1 
MM14 TSMC_28 TSMC_20 TSMC_5 TSMC_5 nch_ulvt_mac l=20n nfin=2 m=1 
XI28 TSMC_15 TSMC_15 TSMC_16 TSMC_5 TSMC_5 TSMC_4 TSMC_3 TSMC_2 
+ S5LLSVTSW8U80_nand3_ulvt_mac_pcell_6 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor3_lvt_mac_pcell_7
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_nor3_lvt_mac_pcell_7 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_9 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_9 TSMC_2 TSMC_10 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_10 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM6 TSMC_8 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_8 TSMC_2 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    vhilo
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_vhilo TSMC_1 TSMC_2 TSMC_3 TSMC_4 
MN3 TSMC_4 TSMC_5 TSMC_6 TSMC_4 nch_svt_mac l=20n nfin=3 m=1 
MN0 TSMC_4 TSMC_6 TSMC_6 TSMC_4 nch_svt_mac l=20n nfin=3 m=1 
MN1 TSMC_4 TSMC_5 TSMC_7 TSMC_4 nch_svt_mac l=20n nfin=3 m=1 
MP7 TSMC_5 TSMC_6 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=3 m=1 
MP2 TSMC_8 TSMC_6 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_5 TSMC_5 TSMC_1 TSMC_1 pch_svt_mac l=20n nfin=3 m=1 
XI16 TSMC_4 TSMC_4 TSMC_8 TSMC_3 TSMC_1 TSMC_1 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI43 TSMC_4 TSMC_4 TSMC_7 TSMC_2 TSMC_1 TSMC_1 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    CKWT_gen
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_CKWT_gen TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 
MM0 TSMC_6 TSMC_10 TSMC_9 TSMC_9 nch_svt_mac l=20n nfin=6 m=7 
MM33 TSMC_4 TSMC_10 TSMC_9 TSMC_9 nch_svt_mac l=20n nfin=6 m=6 
MM51 TSMC_5 TSMC_10 TSMC_9 TSMC_9 nch_svt_mac l=20n nfin=6 m=7 
MM49 TSMC_10 TSMC_2 TSMC_11 TSMC_9 nch_lvt_mac l=16.0n nfin=6 m=8 
MM25 TSMC_10 TSMC_1 TSMC_11 TSMC_9 nch_lvt_mac l=16.0n nfin=6 m=1 
MM53 TSMC_11 TSMC_3 TSMC_9 TSMC_9 nch_lvt_mac l=16.0n nfin=6 m=7 
MM1 TSMC_6 TSMC_10 TSMC_8 TSMC_7 pch_svt_mac l=20n nfin=6 m=7 
MM52 TSMC_5 TSMC_10 TSMC_8 TSMC_7 pch_svt_mac l=20n nfin=6 m=7 
MM34 TSMC_4 TSMC_10 TSMC_8 TSMC_7 pch_svt_mac l=20n nfin=6 m=6 
MM50 TSMC_10 TSMC_3 TSMC_8 TSMC_7 pch_svt_mac l=16.0n nfin=3 m=7 
MM48 TSMC_12 TSMC_2 TSMC_8 TSMC_7 pch_svt_mac l=16.0n nfin=3 m=2 
MM27 TSMC_10 TSMC_1 TSMC_12 TSMC_7 pch_svt_mac l=16.0n nfin=3 m=2 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    ydec_write
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_ydec_write TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 
MM7 TSMC_8 TSMC_2 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=6 m=4 
MM9 TSMC_9 TSMC_1 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=6 m=4 
MM1 TSMC_6 TSMC_9 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=6 m=12 
MM3 TSMC_7 TSMC_8 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=6 m=12 
MM2 TSMC_6 TSMC_9 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=6 m=12 
MM0 TSMC_7 TSMC_8 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=6 m=12 
MM34 TSMC_9 TSMC_1 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=6 m=4 
MM33 TSMC_8 TSMC_2 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=6 m=4 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    ydec_read
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_ydec_read TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM16 TSMC_7 TSMC_9 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=5 m=6 
MM23 TSMC_9 TSMC_6 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=5 m=1 
MM24 TSMC_10 TSMC_6 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=5 m=1 
MM6 TSMC_8 TSMC_10 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=5 m=6 
MM27 TSMC_11 TSMC_2 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=5 m=1 
MM34 TSMC_9 TSMC_11 TSMC_12 TSMC_3 pch_svt_mac l=20n nfin=5 m=2 
MM33 TSMC_10 TSMC_2 TSMC_12 TSMC_3 pch_svt_mac l=20n nfin=5 m=2 
MM17 TSMC_7 TSMC_9 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=5 m=6 
MM25 TSMC_12 TSMC_6 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=5 m=2 
MM5 TSMC_8 TSMC_10 TSMC_4 TSMC_3 pch_svt_mac l=20n nfin=5 m=6 
MM7 TSMC_10 TSMC_2 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=5 m=2 
MM9 TSMC_9 TSMC_11 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=5 m=2 
MM26 TSMC_11 TSMC_2 TSMC_5 TSMC_5 nch_svt_mac l=20n nfin=5 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    rdecb4_wdecb
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_rdecb4_wdecb TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 
MM26 TSMC_12 TSMC_4 TSMC_10 TSMC_9 pch_svt_mac l=20n nfin=3 m=4 
MM1 TSMC_7 TSMC_13 TSMC_10 TSMC_9 pch_svt_mac l=20n nfin=3 m=10 
MM32 TSMC_6 TSMC_14 TSMC_10 TSMC_9 pch_svt_mac l=20n nfin=3 m=10 
MM34 TSMC_5 TSMC_15 TSMC_10 TSMC_9 pch_svt_mac l=20n nfin=3 m=10 
MM2 TSMC_8 TSMC_16 TSMC_10 TSMC_9 pch_svt_mac l=20n nfin=3 m=10 
MM16 TSMC_17 TSMC_3 TSMC_10 TSMC_9 pch_svt_mac l=20n nfin=3 m=4 
MM14 TSMC_13 TSMC_2 TSMC_17 TSMC_9 pch_lvt_mac l=20n nfin=3 m=2 
MM24 TSMC_15 TSMC_2 TSMC_12 TSMC_9 pch_lvt_mac l=20n nfin=3 m=2 
MM25 TSMC_14 TSMC_1 TSMC_12 TSMC_9 pch_lvt_mac l=20n nfin=3 m=2 
MM15 TSMC_16 TSMC_1 TSMC_17 TSMC_9 pch_lvt_mac l=20n nfin=3 m=2 
MM23 TSMC_15 TSMC_2 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
MM22 TSMC_14 TSMC_1 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
MM33 TSMC_6 TSMC_14 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=10 
MM0 TSMC_7 TSMC_13 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=10 
MM19 TSMC_16 TSMC_3 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
MM27 TSMC_15 TSMC_4 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
MM28 TSMC_14 TSMC_4 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
MM18 TSMC_13 TSMC_3 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
MM3 TSMC_8 TSMC_16 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=10 
MM35 TSMC_5 TSMC_15 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=10 
MM13 TSMC_13 TSMC_2 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
MM12 TSMC_16 TSMC_1 TSMC_11 TSMC_11 nch_svt_mac l=20n nfin=3 m=2 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    rdecb4_wdeca
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_rdecb4_wdeca TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
MM55 TSMC_16 TSMC_3 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=8 
MM7 TSMC_17 TSMC_6 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM11 TSMC_18 TSMC_5 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM62 TSMC_9 TSMC_19 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=10 
MM35 TSMC_12 TSMC_20 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=10 
MM29 TSMC_21 TSMC_8 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM27 TSMC_21 TSMC_7 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM4 TSMC_17 TSMC_4 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM23 TSMC_21 TSMC_5 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM28 TSMC_22 TSMC_7 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM22 TSMC_22 TSMC_4 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM54 TSMC_11 TSMC_23 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=10 
MM30 TSMC_22 TSMC_8 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM13 TSMC_18 TSMC_6 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM12 TSMC_18 TSMC_8 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM10 TSMC_17 TSMC_8 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=2 
MM58 TSMC_10 TSMC_24 TSMC_15 TSMC_15 nch_svt_mac l=20n nfin=3 m=10 
MM41 TSMC_20 TSMC_21 TSMC_25 TSMC_15 nch_ulvt_mac l=16.0n nfin=3 m=4 
MM52 TSMC_25 TSMC_2 TSMC_16 TSMC_15 nch_ulvt_mac l=16.0n nfin=3 m=8 
MM16 TSMC_24 TSMC_18 TSMC_25 TSMC_15 nch_ulvt_mac l=16.0n nfin=3 m=4 
MM51 TSMC_25 TSMC_1 TSMC_16 TSMC_15 nch_ulvt_mac l=16.0n nfin=3 m=1 
MM0 TSMC_19 TSMC_17 TSMC_25 TSMC_15 nch_ulvt_mac l=16.0n nfin=3 m=4 
MM32 TSMC_23 TSMC_22 TSMC_25 TSMC_15 nch_ulvt_mac l=16.0n nfin=3 m=4 
MM21 TSMC_25 TSMC_1 TSMC_26 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=1 
MM19 TSMC_20 TSMC_21 TSMC_14 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=2 
MM20 TSMC_26 TSMC_2 TSMC_14 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=1 
MM17 TSMC_24 TSMC_18 TSMC_14 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=2 
MM15 TSMC_19 TSMC_17 TSMC_14 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=2 
MM24 TSMC_25 TSMC_3 TSMC_14 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=1 
MM2 TSMC_27 TSMC_8 TSMC_14 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=6 
MM18 TSMC_23 TSMC_22 TSMC_14 TSMC_13 pch_svt_mac l=16.0n nfin=3 m=2 
MM53 TSMC_11 TSMC_23 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=10 
MM33 TSMC_19 TSMC_3 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=2 
MM8 TSMC_22 TSMC_4 TSMC_28 TSMC_13 pch_ulvt_mac l=20n nfin=3 m=2 
MM9 TSMC_21 TSMC_5 TSMC_28 TSMC_13 pch_ulvt_mac l=20n nfin=3 m=2 
MM25 TSMC_20 TSMC_3 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=2 
MM3 TSMC_17 TSMC_4 TSMC_29 TSMC_13 pch_ulvt_mac l=20n nfin=3 m=2 
MM1 TSMC_29 TSMC_6 TSMC_27 TSMC_13 pch_ulvt_mac l=20n nfin=3 m=4 
MM57 TSMC_10 TSMC_24 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=10 
MM26 TSMC_23 TSMC_3 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=2 
MM34 TSMC_12 TSMC_20 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=10 
MM31 TSMC_24 TSMC_3 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=2 
MM61 TSMC_9 TSMC_19 TSMC_14 TSMC_13 pch_lvt_mac l=20n nfin=3 m=10 
MM14 TSMC_28 TSMC_7 TSMC_27 TSMC_13 pch_ulvt_mac l=20n nfin=3 m=4 
MM6 TSMC_18 TSMC_5 TSMC_29 TSMC_13 pch_ulvt_mac l=20n nfin=3 m=2 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    resetd
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_resetd TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 
MM0 TSMC_11 TSMC_12 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=8 m=1 
MM5 TSMC_4 TSMC_12 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=6 m=6 
MM9 TSMC_1 TSMC_11 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=8 m=6 
MM21 TSMC_7 TSMC_13 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=3 m=1 
MM16 TSMC_12 TSMC_3 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=6 m=4 
MM23 TSMC_6 TSMC_7 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=3 m=2 
MM1 TSMC_11 TSMC_12 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=3 m=2 
MM10 TSMC_1 TSMC_11 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=3 m=12 
MM8 TSMC_4 TSMC_12 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=3 m=12 
MM7 TSMC_12 TSMC_5 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=6 m=4 
XI27 TSMC_4 TSMC_5 TSMC_10 TSMC_10 TSMC_9 TSMC_8 TSMC_13 
+ S5LLSVTSW8U80_nor2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM22 TSMC_7 TSMC_13 TSMC_9 TSMC_8 pch_lvt_mac l=20n nfin=3 m=1 
MM15 TSMC_14 TSMC_3 TSMC_9 TSMC_8 pch_ulvt_mac l=20n nfin=3 m=4 
MM24 TSMC_6 TSMC_7 TSMC_9 TSMC_8 pch_lvt_mac l=20n nfin=3 m=2 
MM6 TSMC_12 TSMC_5 TSMC_14 TSMC_8 pch_ulvt_mac l=20n nfin=3 m=4 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    abufb_lev_x
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_abufb_lev_x TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM9 TSMC_2 TSMC_3 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=6 m=1 
MM5 TSMC_9 TSMC_3 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM6 TSMC_10 TSMC_1 TSMC_11 TSMC_6 pch_svt_mac l=20n nfin=3 m=4 
MM3 TSMC_10 TSMC_4 TSMC_9 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_11 TSMC_5 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=3 m=4 
MM17 TSMC_3 TSMC_10 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=6 m=1 
MM8 TSMC_2 TSMC_3 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=4 m=2 
MM2 TSMC_12 TSMC_4 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=3 m=4 
MM1 TSMC_10 TSMC_5 TSMC_13 TSMC_8 nch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_13 TSMC_3 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=3 m=1 
MM16 TSMC_3 TSMC_10 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=4 m=2 
MM0 TSMC_10 TSMC_1 TSMC_12 TSMC_8 nch_svt_mac l=20n nfin=3 m=4 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    webufb
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_webufb TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 
MM5 TSMC_5 TSMC_3 TSMC_10 TSMC_4 pch_ulvt_mac l=20n nfin=4 m=3 
MP2 TSMC_11 TSMC_2 TSMC_10 TSMC_4 pch_ulvt_mac l=20n nfin=3 m=4 
MM4 TSMC_12 TSMC_1 TSMC_13 TSMC_4 pch_ulvt_mac l=20n nfin=3 m=1 
MP1 TSMC_13 TSMC_7 TSMC_11 TSMC_4 pch_ulvt_mac l=20n nfin=3 m=6 
MP4 TSMC_10 TSMC_14 TSMC_12 TSMC_4 pch_ulvt_mac l=20n nfin=3 m=1 
MTN2 TSMC_15 TSMC_2 TSMC_13 TSMC_6 nch_svt_mac l=20n nfin=3 m=1 
MTN1 TSMC_16 TSMC_1 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=3 m=6 
MTN3 TSMC_6 TSMC_14 TSMC_15 TSMC_6 nch_svt_mac l=20n nfin=3 m=1 
MN0 TSMC_13 TSMC_7 TSMC_16 TSMC_6 nch_svt_mac l=20n nfin=3 m=6 
MM0 TSMC_13 TSMC_3 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=3 m=2 
XI48 TSMC_6 TSMC_6 TSMC_13 TSMC_9 TSMC_5 TSMC_4 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=4 n_nfin=3 n_l=20n p_totalM=4 
+ p_nfin=3 p_l=20n 
XI19 TSMC_6 TSMC_6 TSMC_13 TSMC_14 TSMC_5 TSMC_4 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI20 TSMC_6 TSMC_6 TSMC_14 TSMC_8 TSMC_5 TSMC_4 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=4 n_nfin=3 n_l=20n p_totalM=4 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    abufb_lev_y
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_abufb_lev_y TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM15 TSMC_3 TSMC_9 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=6 m=4 
MM9 TSMC_2 TSMC_10 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=6 m=4 
MM5 TSMC_11 TSMC_10 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=6 m=1 
MM6 TSMC_9 TSMC_1 TSMC_12 TSMC_6 pch_svt_mac l=20n nfin=6 m=2 
MM3 TSMC_9 TSMC_4 TSMC_11 TSMC_6 pch_svt_mac l=20n nfin=6 m=1 
MM4 TSMC_12 TSMC_5 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=6 m=2 
MM17 TSMC_10 TSMC_9 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=6 m=1 
MM8 TSMC_2 TSMC_10 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=6 m=4 
MM14 TSMC_3 TSMC_9 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=6 m=4 
MM2 TSMC_13 TSMC_4 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=6 m=2 
MM1 TSMC_9 TSMC_5 TSMC_14 TSMC_8 nch_svt_mac l=20n nfin=6 m=1 
MM7 TSMC_14 TSMC_10 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=6 m=1 
MM16 TSMC_10 TSMC_9 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=6 m=1 
MM0 TSMC_9 TSMC_1 TSMC_13 TSMC_8 nch_svt_mac l=20n nfin=6 m=2 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    abufb_seg_x
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_abufb_seg_x TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM9 TSMC_2 TSMC_3 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=7 m=1 
MM5 TSMC_9 TSMC_3 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM6 TSMC_10 TSMC_1 TSMC_11 TSMC_6 pch_svt_mac l=20n nfin=3 m=4 
MM3 TSMC_10 TSMC_4 TSMC_9 TSMC_6 pch_svt_mac l=20n nfin=3 m=1 
MM4 TSMC_11 TSMC_5 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=3 m=4 
MM17 TSMC_3 TSMC_10 TSMC_7 TSMC_6 pch_svt_mac l=20n nfin=7 m=1 
MM8 TSMC_2 TSMC_3 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=3 m=2 
MM2 TSMC_12 TSMC_4 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=3 m=4 
MM1 TSMC_10 TSMC_5 TSMC_13 TSMC_8 nch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_13 TSMC_3 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=3 m=1 
MM16 TSMC_3 TSMC_10 TSMC_8 TSMC_8 nch_svt_mac l=20n nfin=3 m=2 
MM0 TSMC_10 TSMC_1 TSMC_12 TSMC_8 nch_svt_mac l=20n nfin=3 m=4 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_ulvt_mac_pcell_8
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_nand2_ulvt_mac_pcell_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    ckp_gen_LS
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_ckp_gen_LS TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 
XI33 TSMC_12 TSMC_13 TSMC_10 TSMC_10 TSMC_9 TSMC_8 TSMC_14 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
MM27 TSMC_15 TSMC_14 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=4 m=1 
MM29 TSMC_2 TSMC_15 TSMC_9 TSMC_8 pch_svt_mac l=20n nfin=4 m=2 
MM19 TSMC_1 TSMC_12 TSMC_16 TSMC_10 nch_svt_mac l=20n nfin=7 m=4 
MM21 TSMC_17 TSMC_1 TSMC_10 TSMC_10 nch_svt_mac l=16.0n nfin=4 m=1 
MM4 TSMC_12 TSMC_4 TSMC_18 TSMC_10 nch_lvt_mac l=20n nfin=8 m=1 
MM30 TSMC_2 TSMC_15 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=4 m=2 
MM20 TSMC_19 TSMC_7 TSMC_17 TSMC_10 nch_svt_mac l=16.0n nfin=4 m=1 
MM22 TSMC_6 TSMC_11 TSMC_10 TSMC_10 nch_svt_mac l=16.0n nfin=8 m=1 
MM28 TSMC_15 TSMC_14 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=4 m=1 
MM3 TSMC_12 TSMC_3 TSMC_18 TSMC_10 nch_lvt_mac l=20n nfin=8 m=1 
MM24 TSMC_6 TSMC_20 TSMC_10 TSMC_10 nch_svt_mac l=16.0n nfin=8 m=1 
MTN3 TSMC_18 TSMC_5 TSMC_21 TSMC_10 nch_lvt_mac l=20n nfin=8 m=1 
MTN2 TSMC_21 TSMC_6 TSMC_10 TSMC_10 nch_lvt_mac l=20n nfin=8 m=1 
MM74 TSMC_16 TSMC_13 TSMC_10 TSMC_10 nch_svt_mac l=20n nfin=7 m=3 
MM17 TSMC_12 TSMC_6 TSMC_9 TSMC_8 pch_ulvt_mac l=20n nfin=8 m=1 
MM11 TSMC_22 TSMC_3 TSMC_9 TSMC_8 pch_ulvt_mac l=16.0n nfin=4 m=1 
MM2 TSMC_23 TSMC_4 TSMC_9 TSMC_8 pch_ulvt_mac l=20n nfin=8 m=1 
MM1 TSMC_12 TSMC_3 TSMC_23 TSMC_8 pch_ulvt_mac l=20n nfin=8 m=1 
MM0 TSMC_12 TSMC_5 TSMC_9 TSMC_8 pch_ulvt_mac l=20n nfin=8 m=1 
MM9 TSMC_19 TSMC_7 TSMC_9 TSMC_8 pch_ulvt_mac l=16.0n nfin=4 m=1 
MM10 TSMC_24 TSMC_4 TSMC_22 TSMC_8 pch_ulvt_mac l=16.0n nfin=4 m=1 
MM13 TSMC_19 TSMC_1 TSMC_9 TSMC_8 pch_ulvt_mac l=16.0n nfin=4 m=1 
M6 TSMC_1 TSMC_13 TSMC_9 TSMC_8 pch_ulvt_mac l=20n nfin=6 m=3 
MM5 TSMC_1 TSMC_12 TSMC_9 TSMC_8 pch_ulvt_mac l=20n nfin=6 m=4 
MM26 TSMC_25 TSMC_11 TSMC_9 TSMC_8 pch_ulvt_mac l=16.0n nfin=8 m=1 
MM25 TSMC_6 TSMC_20 TSMC_25 TSMC_8 pch_ulvt_mac l=16.0n nfin=8 m=1 
MM12 TSMC_24 TSMC_20 TSMC_9 TSMC_8 pch_ulvt_mac l=16.0n nfin=4 m=1 
XI32 TSMC_5 TSMC_6 TSMC_14 TSMC_10 TSMC_10 TSMC_9 TSMC_8 TSMC_13 
+ S5LLSVTSW8U80_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
MM15 TSMC_24 TSMC_4 TSMC_26 TSMC_10 nch_ulvt_mac l=16.0n nfin=4 m=1 
MM16 TSMC_24 TSMC_3 TSMC_26 TSMC_10 nch_ulvt_mac l=16.0n nfin=4 m=1 
MM14 TSMC_26 TSMC_20 TSMC_10 TSMC_10 nch_ulvt_mac l=16.0n nfin=4 m=1 
XI81 TSMC_19 TSMC_24 TSMC_10 TSMC_10 TSMC_9 TSMC_8 TSMC_20 
+ S5LLSVTSW8U80_nand2_ulvt_mac_pcell_8 n_totalM=1 n_nfin=4 n_l=16.0n p_totalM=1 
+ p_nfin=4 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    enbufb_SLP_LS
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_enbufb_SLP_LS TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 
MM69 TSMC_10 TSMC_12 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=4 m=1 
MM81 TSMC_20 TSMC_21 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=6 m=1 
MM68 TSMC_11 TSMC_18 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=8 m=1 
MM64 TSMC_11 TSMC_12 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=8 m=1 
MM74 TSMC_9 TSMC_22 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=7 m=2 
MM76 TSMC_9 TSMC_19 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=2 m=1 
MM77 TSMC_11 TSMC_19 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=2 m=1 
MM78 TSMC_10 TSMC_19 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=2 m=1 
MM79 TSMC_23 TSMC_12 TSMC_20 TSMC_17 nch_svt_mac l=20n nfin=6 m=1 
MM71 TSMC_9 TSMC_12 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=7 m=2 
MM82 TSMC_24 TSMC_8 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=3 m=1 
MM33 TSMC_24 TSMC_1 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=3 m=1 
MM83 TSMC_20 TSMC_19 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=6 m=1 
MM85 TSMC_25 TSMC_14 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=6 m=1 
MM37 TSMC_26 TSMC_14 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=2 m=1 
MM66 TSMC_11 TSMC_22 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=8 m=1 
MM30 TSMC_27 TSMC_13 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=4 m=6 
MTN2 TSMC_12 TSMC_5 TSMC_28 TSMC_17 nch_svt_mac l=20n nfin=8 m=1 
MTN3 TSMC_28 TSMC_26 TSMC_27 TSMC_17 nch_svt_mac l=20n nfin=8 m=1 
MM86 TSMC_22 TSMC_25 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=6 m=2 
MM34 TSMC_26 TSMC_12 TSMC_17 TSMC_17 nch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_29 TSMC_18 TSMC_30 TSMC_15 pch_ulvt_mac l=20n nfin=4 m=4 
MM3 TSMC_30 TSMC_22 TSMC_16 TSMC_15 pch_ulvt_mac l=20n nfin=6 m=4 
MM72 TSMC_9 TSMC_12 TSMC_31 TSMC_15 pch_ulvt_mac l=20n nfin=6 m=2 
M1 TSMC_31 TSMC_22 TSMC_16 TSMC_15 pch_ulvt_mac l=20n nfin=6 m=2 
MM8 TSMC_10 TSMC_12 TSMC_16 TSMC_15 pch_ulvt_mac l=20n nfin=4 m=1 
MM32 TSMC_24 TSMC_1 TSMC_32 TSMC_15 pch_lvt_mac l=20n nfin=3 m=1 
MM9 TSMC_23 TSMC_12 TSMC_16 TSMC_15 pch_ulvt_mac l=20n nfin=12 m=1 
MM12 TSMC_23 TSMC_21 TSMC_33 TSMC_15 pch_ulvt_mac l=20n nfin=12 m=1 
MM75 TSMC_32 TSMC_8 TSMC_16 TSMC_15 pch_lvt_mac l=20n nfin=3 m=1 
MM13 TSMC_33 TSMC_19 TSMC_16 TSMC_15 pch_ulvt_mac l=20n nfin=12 m=1 
MM5 TSMC_11 TSMC_12 TSMC_29 TSMC_15 pch_ulvt_mac l=20n nfin=4 m=4 
MM80 TSMC_25 TSMC_14 TSMC_16 TSMC_15 pch_svt_mac l=20n nfin=6 m=1 
MM36 TSMC_34 TSMC_14 TSMC_16 TSMC_15 pch_svt_mac l=20n nfin=3 m=1 
MM31 TSMC_12 TSMC_13 TSMC_15 TSMC_15 pch_svt_mac l=20n nfin=6 m=1 
MM84 TSMC_22 TSMC_25 TSMC_16 TSMC_15 pch_svt_mac l=20n nfin=6 m=2 
MM35 TSMC_26 TSMC_12 TSMC_34 TSMC_15 pch_svt_mac l=20n nfin=3 m=1 
MP5 TSMC_12 TSMC_2 TSMC_35 TSMC_15 pch_svt_mac l=20n nfin=6 m=1 
MP2 TSMC_36 TSMC_5 TSMC_15 TSMC_15 pch_svt_mac l=20n nfin=8 m=2 
MP4 TSMC_35 TSMC_26 TSMC_15 TSMC_15 pch_svt_mac l=20n nfin=6 m=1 
MP1 TSMC_12 TSMC_24 TSMC_36 TSMC_15 pch_svt_mac l=20n nfin=8 m=2 
MN0 TSMC_12 TSMC_24 TSMC_37 TSMC_17 nch_ulvt_mac l=20n nfin=8 m=2 
MTN1 TSMC_37 TSMC_2 TSMC_27 TSMC_17 nch_ulvt_mac l=20n nfin=8 m=2 
XCKP_GEN TSMC_3 TSMC_4 TSMC_6 TSMC_7 TSMC_23 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_19 S5LLSVTSW8U80_ckp_gen_LS 
XI41 TSMC_17 TSMC_17 TSMC_8 TSMC_21 TSMC_16 TSMC_15 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    cnts2_core_SLP_ls
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_cnts2_core_SLP_ls TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 
XVHILO TSMC_32 TSMC_30 TSMC_31 TSMC_34 S5LLSVTSW8U80_vhilo 
Xckwt_gen<0> TSMC_13 TSMC_15 TSMC_20 TSMC_21 TSMC_23 TSMC_24 TSMC_32 TSMC_32 
+ TSMC_34 S5LLSVTSW8U80_CKWT_gen 
Xckwt_gen<1> TSMC_13 TSMC_15 TSMC_20 TSMC_22 TSMC_25 TSMC_26 TSMC_32 TSMC_32 
+ TSMC_34 S5LLSVTSW8U80_CKWT_gen 
XYDEC_WRITE<0> TSMC_10 TSMC_9 TSMC_32 TSMC_33 TSMC_34 TSMC_58 TSMC_59 
+ S5LLSVTSW8U80_ydec_write 
XYDEC_WRITE<1> TSMC_10 TSMC_9 TSMC_32 TSMC_33 TSMC_34 TSMC_60 TSMC_61 
+ S5LLSVTSW8U80_ydec_write 
XYDEC_READ<0> TSMC_10 TSMC_9 TSMC_32 TSMC_33 TSMC_34 TSMC_52 TSMC_54 
+ TSMC_55 S5LLSVTSW8U80_ydec_read 
XYDEC_READ<1> TSMC_10 TSMC_9 TSMC_32 TSMC_33 TSMC_34 TSMC_52 TSMC_56 
+ TSMC_57 S5LLSVTSW8U80_ydec_read 
XRDECB4_WDECB TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_32 TSMC_33 TSMC_34 S5LLSVTSW8U80_rdecb4_wdecb 
XRDECB4_WDECC TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_47 TSMC_48 TSMC_49 
+ TSMC_50 TSMC_32 TSMC_33 TSMC_34 S5LLSVTSW8U80_rdecb4_wdecb 
XRDECB4_WDECA<0> TSMC_13 TSMC_15 TSMC_19 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_75 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_rdecb4_wdeca 
XRDECB4_WDECA<1> TSMC_13 TSMC_15 TSMC_19 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_76 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_rdecb4_wdeca 
XRESETD TSMC_12 TSMC_13 TSMC_14 TSMC_77 TSMC_16 TSMC_78 TSMC_79 TSMC_32 TSMC_33 
+ TSMC_34 S5LLSVTSW8U80_resetd 
XABUFB_DECB<0> TSMC_5 TSMC_63 TSMC_64 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_lev_x 
XABUFB_DECB<1> TSMC_6 TSMC_65 TSMC_66 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_lev_x 
XABUFB_DECC<0> TSMC_7 TSMC_67 TSMC_68 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_lev_x 
XABUFB_DECC<1> TSMC_8 TSMC_69 TSMC_70 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_lev_x 
XWEBUFB TSMC_12 TSMC_77 TSMC_17 TSMC_32 TSMC_33 TSMC_34 TSMC_51 TSMC_52 TSMC_53 
+ S5LLSVTSW8U80_webufb 
XABUFB_YDECW TSMC_1 TSMC_9 TSMC_10 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_lev_y 
XABUFB_DECA<0> TSMC_2 TSMC_72 TSMC_71 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_seg_x 
XABUFB_DECA<1> TSMC_3 TSMC_74 TSMC_73 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_seg_x 
XABUFB_DECA<2> TSMC_4 TSMC_76 TSMC_75 TSMC_12 TSMC_77 TSMC_32 TSMC_33 TSMC_34 
+ S5LLSVTSW8U80_abufb_seg_x 
XENBUFB TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_77 TSMC_15 TSMC_16 TSMC_17 TSMC_19 
+ TSMC_18 TSMC_20 TSMC_27 TSMC_28 TSMC_29 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_53 TSMC_62 S5LLSVTSW8U80_enbufb_SLP_LS 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    xdel_sae_slp_MUX1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_xdel_sae_slp_MUX1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 
MM110 TSMC_28 TSMC_29 TSMC_19 TSMC_18 pch_svt_mac l=20n nfin=6 m=1 
MM109 TSMC_10 TSMC_30 TSMC_18 TSMC_18 pch_svt_mac l=16.0n nfin=6 m=2 
MM105 TSMC_8 TSMC_31 TSMC_18 TSMC_18 pch_svt_mac l=16.0n nfin=6 m=2 
MM103 TSMC_9 TSMC_30 TSMC_18 TSMC_18 pch_svt_mac l=16.0n nfin=6 m=2 
MM21 TSMC_30 TSMC_32 TSMC_19 TSMC_18 pch_lvt_mac l=16.0n nfin=7 m=2 
MM88 TSMC_33 TSMC_5 TSMC_34 TSMC_18 pch_lvt_mac l=16.0n nfin=6 m=1 
MM18 TSMC_35 TSMC_3 TSMC_19 TSMC_18 pch_lvt_mac l=16.0n nfin=6 m=1 
MM17 TSMC_33 TSMC_2 TSMC_35 TSMC_18 pch_lvt_mac l=16.0n nfin=6 m=1 
MM86 TSMC_33 TSMC_36 TSMC_19 TSMC_18 pch_lvt_mac l=16.0n nfin=6 m=1 
MM72 TSMC_32 TSMC_37 TSMC_18 TSMC_18 pch_svt_mac l=16.0n nfin=6 m=1 
MM73 TSMC_32 TSMC_38 TSMC_18 TSMC_18 pch_svt_mac l=16.0n nfin=6 m=1 
MM71 TSMC_39 TSMC_13 TSMC_19 TSMC_18 pch_svt_mac l=20n nfin=3 m=1 
MM75 TSMC_32 TSMC_40 TSMC_18 TSMC_18 pch_svt_mac l=16.0n nfin=6 m=1 
MM95 TSMC_7 TSMC_31 TSMC_18 TSMC_18 pch_svt_mac l=16.0n nfin=6 m=2 
MM33 TSMC_8 TSMC_31 TSMC_18 TSMC_18 pch_svt_mac l=20n nfin=6 m=6 
MM92 TSMC_34 TSMC_1 TSMC_19 TSMC_18 pch_lvt_mac l=16.0n nfin=6 m=1 
MM23 TSMC_31 TSMC_32 TSMC_19 TSMC_18 pch_lvt_mac l=16.0n nfin=7 m=2 
MM37 TSMC_9 TSMC_30 TSMC_18 TSMC_18 pch_svt_mac l=20n nfin=6 m=6 
MM12 TSMC_7 TSMC_31 TSMC_18 TSMC_18 pch_svt_mac l=20n nfin=6 m=6 
MM35 TSMC_10 TSMC_30 TSMC_18 TSMC_18 pch_svt_mac l=20n nfin=6 m=6 
MM116 TSMC_41 TSMC_37 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=2 m=1 
MM113 TSMC_42 TSMC_37 TSMC_41 TSMC_20 nch_svt_mac l=20n nfin=2 m=1 
MM106 TSMC_37 TSMC_17 TSMC_43 TSMC_20 nch_svt_mac l=16.0n nfin=3 m=3 
MM104 TSMC_43 TSMC_44 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=3 m=2 
MM96 TSMC_30 TSMC_32 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=6 m=2 
MM94 TSMC_45 TSMC_33 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=4 m=1 
MM91 TSMC_16 TSMC_33 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=4 m=1 
MM90 TSMC_16 TSMC_21 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=4 m=1 
MM89 TSMC_14 TSMC_46 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=3 m=1 
MM87 TSMC_47 TSMC_5 TSMC_20 TSMC_20 nch_lvt_mac l=16.0n nfin=9 m=1 
MM15 TSMC_33 TSMC_2 TSMC_48 TSMC_20 nch_lvt_mac l=16.0n nfin=9 m=1 
MM16 TSMC_33 TSMC_3 TSMC_48 TSMC_20 nch_lvt_mac l=16.0n nfin=9 m=1 
MM98 TSMC_7 TSMC_31 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=9 m=4 
MM100 TSMC_8 TSMC_31 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=9 m=4 
MM74 TSMC_14 TSMC_45 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=2 m=3 
MM78 TSMC_40 TSMC_1 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=3 m=1 
MM79 TSMC_40 TSMC_21 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=3 m=1 
MM93 TSMC_45 TSMC_22 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=4 m=1 
MM101 TSMC_10 TSMC_30 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=9 m=4 
MM159 TSMC_31 TSMC_23 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=2 m=2 
MM162 TSMC_30 TSMC_23 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=2 m=2 
MM102 TSMC_37 TSMC_14 TSMC_43 TSMC_20 nch_svt_mac l=16.0n nfin=3 m=2 
MM97 TSMC_31 TSMC_32 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=6 m=2 
MM14 TSMC_48 TSMC_36 TSMC_47 TSMC_20 nch_lvt_mac l=16.0n nfin=9 m=1 
MM111 TSMC_49 TSMC_42 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=2 m=1 
MM61 TSMC_50 TSMC_49 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=2 m=3 
MM60 TSMC_38 TSMC_32 TSMC_50 TSMC_20 nch_svt_mac l=20n nfin=2 m=3 
MM80 TSMC_51 TSMC_13 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=3 m=1 
MM99 TSMC_9 TSMC_30 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=9 m=4 
MM77 TSMC_40 TSMC_23 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=3 m=1 
MM57 TSMC_38 TSMC_11 TSMC_50 TSMC_20 nch_svt_mac l=20n nfin=2 m=3 
MM34 TSMC_10 TSMC_30 TSMC_20 TSMC_20 nch_lvt_mac l=20n nfin=6 m=6 
MM36 TSMC_9 TSMC_30 TSMC_20 TSMC_20 nch_lvt_mac l=20n nfin=6 m=6 
MM232 TSMC_6 TSMC_51 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=3 m=4 
MM11 TSMC_7 TSMC_31 TSMC_20 TSMC_20 nch_lvt_mac l=20n nfin=6 m=6 
MM47 TSMC_46 TSMC_33 TSMC_20 TSMC_20 nch_svt_mac l=16.0n nfin=3 m=1 
MM108 TSMC_44 TSMC_29 TSMC_20 TSMC_20 nch_svt_mac l=20n nfin=3 m=1 
MM63 TSMC_37 TSMC_33 TSMC_20 TSMC_20 nch_lvt_mac l=16.0n nfin=2 m=3 
MM32 TSMC_8 TSMC_31 TSMC_20 TSMC_20 nch_lvt_mac l=20n nfin=6 m=6 
MM107 TSMC_47 TSMC_1 TSMC_20 TSMC_20 nch_lvt_mac l=16.0n nfin=9 m=1 
Xresetd_tsel TSMC_2 TSMC_36 TSMC_13 TSMC_18 TSMC_19 TSMC_20 TSMC_24 TSMC_25 
+ S5LLSVTSW8U80_RESETD_RTSEL 
XI128 TSMC_37 TSMC_52 TSMC_20 TSMC_20 TSMC_39 TSMC_18 TSMC_51 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
Xresetd_rtsel TSMC_37 TSMC_52 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_26 TSMC_27 
+ S5LLSVTSW8U80_RESETD_WTSEL 
XI139 TSMC_20 TSMC_20 TSMC_17 TSMC_53 TSMC_19 TSMC_18 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI141 TSMC_20 TSMC_20 TSMC_4 TSMC_54 TSMC_28 TSMC_18 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI154 TSMC_54 TSMC_46 TSMC_17 TSMC_20 TSMC_20 TSMC_28 TSMC_18 TSMC_44 
+ S5LLSVTSW8U80_nand3_lvt_mac_pcell_2 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI164 TSMC_24 TSMC_25 TSMC_17 TSMC_20 TSMC_20 TSMC_19 TSMC_18 TSMC_29 
+ S5LLSVTSW8U80_nor3_lvt_mac_pcell_7 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
MM3 TSMC_49 TSMC_42 TSMC_19 TSMC_18 pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_55 TSMC_37 TSMC_19 TSMC_18 pch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_42 TSMC_37 TSMC_55 TSMC_18 pch_svt_mac l=20n nfin=2 m=1 
MM62 TSMC_38 TSMC_49 TSMC_19 TSMC_18 pch_svt_mac l=20n nfin=3 m=1 
MM22 TSMC_6 TSMC_51 TSMC_19 TSMC_18 pch_svt_mac l=20n nfin=2 m=4 
MM6 TSMC_15 TSMC_33 TSMC_19 TSMC_18 pch_ulvt_mac l=20n nfin=5 m=2 
MM31 TSMC_56 TSMC_17 TSMC_57 TSMC_18 pch_lvt_mac l=16.0n nfin=3 m=3 
MM59 TSMC_58 TSMC_32 TSMC_19 TSMC_18 pch_ulvt_mac l=20n nfin=3 m=1 
MM27 TSMC_37 TSMC_14 TSMC_56 TSMC_18 pch_lvt_mac l=16.0n nfin=4 m=2 
MM26 TSMC_37 TSMC_44 TSMC_57 TSMC_18 pch_lvt_mac l=16.0n nfin=4 m=2 
MM19 TSMC_45 TSMC_33 TSMC_59 TSMC_18 pch_ulvt_mac l=16.0n nfin=6 m=1 
MM10 TSMC_16 TSMC_33 TSMC_60 TSMC_18 pch_ulvt_mac l=16.0n nfin=6 m=2 
MM9 TSMC_60 TSMC_21 TSMC_19 TSMC_18 pch_ulvt_mac l=16.0n nfin=6 m=2 
MM13 TSMC_59 TSMC_22 TSMC_19 TSMC_18 pch_ulvt_mac l=16.0n nfin=6 m=1 
MM2 TSMC_40 TSMC_21 TSMC_61 TSMC_18 pch_ulvt_mac l=20n nfin=6 m=1 
MM0 TSMC_62 TSMC_23 TSMC_19 TSMC_18 pch_ulvt_mac l=20n nfin=6 m=1 
MM1 TSMC_61 TSMC_1 TSMC_62 TSMC_18 pch_ulvt_mac l=20n nfin=6 m=1 
MM39 TSMC_14 TSMC_46 TSMC_19 TSMC_18 pch_ulvt_mac l=16.0n nfin=3 m=4 
MM25 TSMC_57 TSMC_33 TSMC_19 TSMC_18 pch_lvt_mac l=16.0n nfin=3 m=3 
MM58 TSMC_38 TSMC_11 TSMC_58 TSMC_18 pch_ulvt_mac l=20n nfin=3 m=1 
MM50 TSMC_46 TSMC_33 TSMC_19 TSMC_18 pch_ulvt_mac l=16.0n nfin=3 m=1 
MM117 TSMC_15 TSMC_33 TSMC_20 TSMC_20 nch_ulvt_mac l=20n nfin=5 m=2 
MM82 TSMC_63 TSMC_38 TSMC_64 TSMC_20 nch_ulvt_mac l=16.0n nfin=10 m=1 
MM83 TSMC_64 TSMC_40 TSMC_20 TSMC_20 nch_ulvt_mac l=16.0n nfin=10 m=1 
MM81 TSMC_32 TSMC_37 TSMC_63 TSMC_20 nch_ulvt_mac l=16.0n nfin=10 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    lctrl_l_core_slp_MUX1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_lctrl_l_core_slp_MUX1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
MM149 TSMC_34 TSMC_35 TSMC_27 TSMC_26 pch_ulvt_mac l=20n nfin=6 m=4 
MM151 TSMC_36 TSMC_35 TSMC_27 TSMC_26 pch_ulvt_mac l=20n nfin=6 m=4 
MM90 TSMC_18 TSMC_36 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=6 m=5 
MM107 TSMC_35 TSMC_2 TSMC_37 TSMC_28 nch_ulvt_mac l=20n nfin=6 m=1 
MM150 TSMC_36 TSMC_35 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=3 m=4 
MM159 TSMC_34 TSMC_33 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=2 m=1 
MM152 TSMC_37 TSMC_6 TSMC_28 TSMC_28 nch_ulvt_mac l=20n nfin=6 m=4 
MM41 TSMC_16 TSMC_34 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=6 m=5 
MM30 TSMC_17 TSMC_34 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=6 m=5 
MM36 TSMC_35 TSMC_4 TSMC_37 TSMC_28 nch_ulvt_mac l=20n nfin=6 m=4 
MM88 TSMC_19 TSMC_36 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=6 m=5 
MM162 TSMC_36 TSMC_33 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=2 m=1 
MM148 TSMC_34 TSMC_35 TSMC_28 TSMC_28 nch_svt_mac l=20n nfin=3 m=4 
MM91 TSMC_18 TSMC_36 TSMC_26 TSMC_26 pch_svt_mac l=20n nfin=6 m=5 
MM89 TSMC_19 TSMC_36 TSMC_26 TSMC_26 pch_svt_mac l=20n nfin=6 m=5 
MM161 TSMC_35 TSMC_6 TSMC_26 TSMC_26 pch_svt_mac l=20n nfin=6 m=1 
MM108 TSMC_38 TSMC_4 TSMC_26 TSMC_26 pch_svt_mac l=20n nfin=6 m=1 
MM40 TSMC_16 TSMC_34 TSMC_26 TSMC_26 pch_svt_mac l=20n nfin=6 m=5 
MM37 TSMC_35 TSMC_2 TSMC_38 TSMC_26 pch_svt_mac l=20n nfin=6 m=1 
MM35 TSMC_17 TSMC_34 TSMC_26 TSMC_26 pch_svt_mac l=20n nfin=6 m=5 
Xxdel_sae TSMC_1 TSMC_2 TSMC_4 TSMC_5 TSMC_7 TSMC_8 TSMC_11 TSMC_12 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_33 TSMC_9 TSMC_10 
+ TSMC_31 TSMC_32 S5LLSVTSW8U80_xdel_sae_slp_MUX1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    lctrl_l_slp_MUX1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_lctrl_l_slp_MUX1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
XLCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ S5LLSVTSW8U80_lctrl_l_core_slp_MUX1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    BIT1A_L20
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_BIT1A_L20 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 
XIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_18 TSMC_19 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_16 
+ TSMC_16 TSMC_17 S5LLSVTSW8U80_BIT1A_CORE_L20 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    CNTS1_SLP
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_CNTS1_SLP TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
XI209<0> TSMC_64 TSMC_64 TSMC_41 TSMC_86 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI209<1> TSMC_64 TSMC_64 TSMC_42 TSMC_87 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI236 TSMC_64 TSMC_64 TSMC_48 TSMC_49 TSMC_88 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI211<0> TSMC_64 TSMC_64 TSMC_84 TSMC_89 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI211<1> TSMC_64 TSMC_64 TSMC_85 TSMC_90 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI212<0> TSMC_64 TSMC_64 TSMC_86 TSMC_91 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI212<1> TSMC_64 TSMC_64 TSMC_87 TSMC_92 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI214<0> TSMC_64 TSMC_64 TSMC_89 TSMC_93 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI214<1> TSMC_64 TSMC_64 TSMC_90 TSMC_94 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI220 TSMC_64 TSMC_64 TSMC_61 TSMC_95 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI241<0> TSMC_64 TSMC_64 TSMC_15 TSMC_96 TSMC_97 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI241<1> TSMC_64 TSMC_64 TSMC_16 TSMC_98 TSMC_97 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI221 TSMC_64 TSMC_64 TSMC_95 TSMC_99 TSMC_63 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI251<0> TSMC_64 TSMC_64 TSMC_96 TSMC_17 TSMC_97 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI251<1> TSMC_64 TSMC_64 TSMC_98 TSMC_18 TSMC_97 TSMC_62 
+ S5LLSVTSW8U80_inv_lvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI247 TSMC_48 TSMC_13 TSMC_64 TSMC_64 TSMC_62 TSMC_62 TSMC_14 
+ S5LLSVTSW8U80_nor2_lvt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
MM12 TSMC_88 TSMC_48 TSMC_62 TSMC_62 pch_svt_mac l=20n nfin=2 m=1 
MM38 TSMC_97 TSMC_48 TSMC_62 TSMC_62 pch_svt_mac l=20n nfin=2 m=1 
XCNT TSMC_57 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_100 TSMC_101 
+ TSMC_9 TSMC_102 TSMC_10 TSMC_103 TSMC_11 TSMC_11 TSMC_8 TSMC_19 
+ TSMC_104 TSMC_105 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_38 TSMC_39 TSMC_40 TSMC_56 TSMC_57 TSMC_62 TSMC_63 TSMC_64 
+ TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 
+ TSMC_82 TSMC_83 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 TSMC_113 TSMC_12 S5LLSVTSW8U80_cnts2_core_SLP_ls 
MM6 TSMC_67 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
MM0 TSMC_23 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=2 m=2 
MM2 TSMC_25 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=2 m=2 
MM1 TSMC_24 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=2 m=2 
MM4 TSMC_66 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_65 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
MM8 TSMC_22 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=2 m=2 
MM10 TSMC_72 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
MM11 TSMC_71 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
MM5 TSMC_68 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
MM9 TSMC_70 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_69 TSMC_12 TSMC_64 TSMC_64 nch_svt_mac l=20n nfin=3 m=1 
XLCTRL TSMC_8 TSMC_10 TSMC_103 TSMC_11 TSMC_11 TSMC_19 TSMC_104 TSMC_40 TSMC_91 
+ TSMC_92 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_99 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_82 TSMC_83 TSMC_93 TSMC_94 TSMC_12 
+ S5LLSVTSW8U80_lctrl_l_slp_MUX1 
XI249 TSMC_14 TSMC_54 TSMC_64 TSMC_64 TSMC_62 TSMC_62 TSMC_55 
+ S5LLSVTSW8U80_nand2_lvt_mac_pcell_4 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    DIOA
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_DIOA TSMC_1 TSMC_2 TSMC_3 
MM0 TSMC_1 TSMC_2 TSMC_1 TSMC_3 nch_svt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: n16ff_uhd1prf_sb_leafcell
* Cell Name:    IOEDGE_L_MUX1
* View Name:    schematic
************************************************************************

.SUBCKT S5LLSVTSW8U80_IOEDGE_L_MUX1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
MM36 TSMC_7 TSMC_2 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=3 m=1 
MM0 TSMC_3 TSMC_8 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=2 m=10 
MM117 TSMC_8 TSMC_7 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=2 m=2 
MM115 TSMC_7 TSMC_1 TSMC_6 TSMC_6 nch_svt_mac l=20n nfin=3 m=1 
MM28 TSMC_9 TSMC_2 TSMC_5 TSMC_4 pch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_3 TSMC_8 TSMC_5 TSMC_4 pch_svt_mac l=20n nfin=2 m=10 
MM118 TSMC_8 TSMC_7 TSMC_5 TSMC_4 pch_svt_mac l=20n nfin=2 m=2 
MM116 TSMC_7 TSMC_1 TSMC_9 TSMC_4 pch_svt_mac l=20n nfin=3 m=1 
.ENDS

.SUBCKT S5LLSVTSW8U80_DIOBIT TSMC_1 TSMC_2 
XD1 TSMC_2 TSMC_1 ndio_mac nfin=2 l=2e-07 m=1 
.ENDS

.SUBCKT ndio_mac PLUS MINUS 
.ENDS



**** End of leaf cells

.SUBCKT S5LLSVTSW8U80_MCB_1X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 
XMCB_0 TSMC_1 TSMC_3 TSMC_5 TSMC_7 TSMC_8 TSMC_9 
+ S5LLSVTSW8U80_MCB_D0907 
XMCB_1 TSMC_2 TSMC_4 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ S5LLSVTSW8U80_MCB_D0907 
.ENDS

.SUBCKT S5LLSVTSW8U80_MCB_2X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 
XMCB_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ S5LLSVTSW8U80_MCB_1X2 
XMCB_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_10 
+ S5LLSVTSW8U80_MCB_1X2 
.ENDS

.SUBCKT S5LLSVTSW8U80_MCB_ARR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
XMCB_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 S5LLSVTSW8U80_MCB_2X2 
XMCB_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_11 
+ TSMC_12 S5LLSVTSW8U80_MCB_2X2 
XMCB_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_13 
+ TSMC_14 S5LLSVTSW8U80_MCB_2X2 
XMCB_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_15 
+ TSMC_16 S5LLSVTSW8U80_MCB_2X2 
.ENDS

.SUBCKT S5LLSVTSW8U80_TKBL_ARR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XTKBL_ON_CELL_0 TSMC_1 TSMC_2 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_13 
+ TSMC_12 S5LLSVTSW8U80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_1 TSMC_1 TSMC_2 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_11 
+ TSMC_10 S5LLSVTSW8U80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_2 TSMC_1 TSMC_2 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_9 TSMC_8 
+ S5LLSVTSW8U80_MCB_D0907_ONCELL 
XTKBL_ON_CELL_3 TSMC_1 TSMC_2 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_7 TSMC_6 
+ S5LLSVTSW8U80_MCB_D0907_ONCELL 
.ENDS

.SUBCKT S5LLSVTSW8U80_MIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
XBIT1A TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_11 TSMC_12 
+ TSMC_9 TSMC_10 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ S5LLSVTSW8U80_BIT1A_L20 
.ENDS

.SUBCKT TS5N16FFCLLSVTA8X128M1SW A[0] A[1] A[2] BWEB[0] BWEB[1] BWEB[2] BWEB[3] 
+ BWEB[4] BWEB[5] BWEB[6] BWEB[7] BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12] 
+ BWEB[13] BWEB[14] BWEB[15] BWEB[16] BWEB[17] BWEB[18] BWEB[19] BWEB[20] 
+ BWEB[21] BWEB[22] BWEB[23] BWEB[24] BWEB[25] BWEB[26] BWEB[27] BWEB[28] 
+ BWEB[29] BWEB[30] BWEB[31] BWEB[32] BWEB[33] BWEB[34] BWEB[35] BWEB[36] 
+ BWEB[37] BWEB[38] BWEB[39] BWEB[40] BWEB[41] BWEB[42] BWEB[43] BWEB[44] 
+ BWEB[45] BWEB[46] BWEB[47] BWEB[48] BWEB[49] BWEB[50] BWEB[51] BWEB[52] 
+ BWEB[53] BWEB[54] BWEB[55] BWEB[56] BWEB[57] BWEB[58] BWEB[59] BWEB[60] 
+ BWEB[61] BWEB[62] BWEB[63] BWEB[64] BWEB[65] BWEB[66] BWEB[67] BWEB[68] 
+ BWEB[69] BWEB[70] BWEB[71] BWEB[72] BWEB[73] BWEB[74] BWEB[75] BWEB[76] 
+ BWEB[77] BWEB[78] BWEB[79] BWEB[80] BWEB[81] BWEB[82] BWEB[83] BWEB[84] 
+ BWEB[85] BWEB[86] BWEB[87] BWEB[88] BWEB[89] BWEB[90] BWEB[91] BWEB[92] 
+ BWEB[93] BWEB[94] BWEB[95] BWEB[96] BWEB[97] BWEB[98] BWEB[99] BWEB[100] 
+ BWEB[101] BWEB[102] BWEB[103] BWEB[104] BWEB[105] BWEB[106] BWEB[107] 
+ BWEB[108] BWEB[109] BWEB[110] BWEB[111] BWEB[112] BWEB[113] BWEB[114] 
+ BWEB[115] BWEB[116] BWEB[117] BWEB[118] BWEB[119] BWEB[120] BWEB[121] 
+ BWEB[122] BWEB[123] BWEB[124] BWEB[125] BWEB[126] BWEB[127] D[0] D[1] D[2] 
+ D[3] D[4] D[5] D[6] D[7] D[8] D[9] D[10] D[11] D[12] D[13] D[14] D[15] D[16] 
+ D[17] D[18] D[19] D[20] D[21] D[22] D[23] D[24] D[25] D[26] D[27] D[28] D[29] 
+ D[30] D[31] D[32] D[33] D[34] D[35] D[36] D[37] D[38] D[39] D[40] D[41] D[42] 
+ D[43] D[44] D[45] D[46] D[47] D[48] D[49] D[50] D[51] D[52] D[53] D[54] D[55] 
+ D[56] D[57] D[58] D[59] D[60] D[61] D[62] D[63] D[64] D[65] D[66] D[67] D[68] 
+ D[69] D[70] D[71] D[72] D[73] D[74] D[75] D[76] D[77] D[78] D[79] D[80] D[81] 
+ D[82] D[83] D[84] D[85] D[86] D[87] D[88] D[89] D[90] D[91] D[92] D[93] D[94] 
+ D[95] D[96] D[97] D[98] D[99] D[100] D[101] D[102] D[103] D[104] D[105] 
+ D[106] D[107] D[108] D[109] D[110] D[111] D[112] D[113] D[114] D[115] D[116] 
+ D[117] D[118] D[119] D[120] D[121] D[122] D[123] D[124] D[125] D[126] D[127] 
+ Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] Q[11] Q[12] Q[13] 
+ Q[14] Q[15] Q[16] Q[17] Q[18] Q[19] Q[20] Q[21] Q[22] Q[23] Q[24] Q[25] Q[26] 
+ Q[27] Q[28] Q[29] Q[30] Q[31] Q[32] Q[33] Q[34] Q[35] Q[36] Q[37] Q[38] Q[39] 
+ Q[40] Q[41] Q[42] Q[43] Q[44] Q[45] Q[46] Q[47] Q[48] Q[49] Q[50] Q[51] Q[52] 
+ Q[53] Q[54] Q[55] Q[56] Q[57] Q[58] Q[59] Q[60] Q[61] Q[62] Q[63] Q[64] Q[65] 
+ Q[66] Q[67] Q[68] Q[69] Q[70] Q[71] Q[72] Q[73] Q[74] Q[75] Q[76] Q[77] Q[78] 
+ Q[79] Q[80] Q[81] Q[82] Q[83] Q[84] Q[85] Q[86] Q[87] Q[88] Q[89] Q[90] Q[91] 
+ Q[92] Q[93] Q[94] Q[95] Q[96] Q[97] Q[98] Q[99] Q[100] Q[101] Q[102] Q[103] 
+ Q[104] Q[105] Q[106] Q[107] Q[108] Q[109] Q[110] Q[111] Q[112] Q[113] Q[114] 
+ Q[115] Q[116] Q[117] Q[118] Q[119] Q[120] Q[121] Q[122] Q[123] Q[124] Q[125] 
+ Q[126] Q[127] RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] VDD VSS WEB CEB CLK 
XMCB8_L_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_1 TSMC_13 TSMC_14 TSMC_15 TSMC_16 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_2 TSMC_17 TSMC_18 TSMC_19 TSMC_20 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_3 TSMC_21 TSMC_22 TSMC_23 TSMC_24 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_4 TSMC_25 TSMC_26 TSMC_27 TSMC_28 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_5 TSMC_29 TSMC_30 TSMC_31 TSMC_32 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_6 TSMC_33 TSMC_34 TSMC_35 TSMC_36 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_7 TSMC_37 TSMC_38 TSMC_39 TSMC_40 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_8 TSMC_41 TSMC_42 TSMC_43 TSMC_44 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_9 TSMC_45 TSMC_46 TSMC_47 TSMC_48 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_10 TSMC_49 TSMC_50 TSMC_51 TSMC_52 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_11 TSMC_53 TSMC_54 TSMC_55 TSMC_56 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_12 TSMC_57 TSMC_58 TSMC_59 TSMC_60 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_13 TSMC_61 TSMC_62 TSMC_63 TSMC_64 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_14 TSMC_65 TSMC_66 TSMC_67 TSMC_68 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_15 TSMC_69 TSMC_70 TSMC_71 TSMC_72 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_16 TSMC_73 TSMC_74 TSMC_75 TSMC_76 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_17 TSMC_77 TSMC_78 TSMC_79 TSMC_80 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_18 TSMC_81 TSMC_82 TSMC_83 TSMC_84 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_19 TSMC_85 TSMC_86 TSMC_87 TSMC_88 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_20 TSMC_89 TSMC_90 TSMC_91 TSMC_92 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_21 TSMC_93 TSMC_94 TSMC_95 TSMC_96 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_22 TSMC_97 TSMC_98 TSMC_99 TSMC_100 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_23 TSMC_101 TSMC_102 TSMC_103 TSMC_104 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_24 TSMC_105 TSMC_106 TSMC_107 TSMC_108 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_25 TSMC_109 TSMC_110 TSMC_111 TSMC_112 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_26 TSMC_113 TSMC_114 TSMC_115 TSMC_116 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_27 TSMC_117 TSMC_118 TSMC_119 TSMC_120 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_28 TSMC_121 TSMC_122 TSMC_123 TSMC_124 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_29 TSMC_125 TSMC_126 TSMC_127 TSMC_128 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_30 TSMC_129 TSMC_130 TSMC_131 TSMC_132 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_L_31 TSMC_133 TSMC_134 TSMC_135 TSMC_136 VDD VDD VDD VSS TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_32 TSMC_137 TSMC_138 TSMC_139 TSMC_140 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_33 TSMC_149 TSMC_150 TSMC_151 TSMC_152 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_34 TSMC_153 TSMC_154 TSMC_155 TSMC_156 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_35 TSMC_157 TSMC_158 TSMC_159 TSMC_160 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_36 TSMC_161 TSMC_162 TSMC_163 TSMC_164 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_37 TSMC_165 TSMC_166 TSMC_167 TSMC_168 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_38 TSMC_169 TSMC_170 TSMC_171 TSMC_172 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_39 TSMC_173 TSMC_174 TSMC_175 TSMC_176 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_40 TSMC_177 TSMC_178 TSMC_179 TSMC_180 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_41 TSMC_181 TSMC_182 TSMC_183 TSMC_184 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_42 TSMC_185 TSMC_186 TSMC_187 TSMC_188 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_43 TSMC_189 TSMC_190 TSMC_191 TSMC_192 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_44 TSMC_193 TSMC_194 TSMC_195 TSMC_196 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_45 TSMC_197 TSMC_198 TSMC_199 TSMC_200 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_46 TSMC_201 TSMC_202 TSMC_203 TSMC_204 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_47 TSMC_205 TSMC_206 TSMC_207 TSMC_208 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_48 TSMC_209 TSMC_210 TSMC_211 TSMC_212 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_49 TSMC_213 TSMC_214 TSMC_215 TSMC_216 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_50 TSMC_217 TSMC_218 TSMC_219 TSMC_220 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_51 TSMC_221 TSMC_222 TSMC_223 TSMC_224 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_52 TSMC_225 TSMC_226 TSMC_227 TSMC_228 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_53 TSMC_229 TSMC_230 TSMC_231 TSMC_232 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_54 TSMC_233 TSMC_234 TSMC_235 TSMC_236 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_55 TSMC_237 TSMC_238 TSMC_239 TSMC_240 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_56 TSMC_241 TSMC_242 TSMC_243 TSMC_244 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_57 TSMC_245 TSMC_246 TSMC_247 TSMC_248 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_58 TSMC_249 TSMC_250 TSMC_251 TSMC_252 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_59 TSMC_253 TSMC_254 TSMC_255 TSMC_256 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_60 TSMC_257 TSMC_258 TSMC_259 TSMC_260 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_61 TSMC_261 TSMC_262 TSMC_263 TSMC_264 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_62 TSMC_265 TSMC_266 TSMC_267 TSMC_268 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XMCB8_R_63 TSMC_269 TSMC_270 TSMC_271 TSMC_272 VDD VDD VDD VSS TSMC_141 
+ TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_MCB_ARR 
XWLDVX1_L0 VDD VSS TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ S5LLSVTSW8U80_WLDRV4X1 
XWLDVX1_L1 VDD VSS TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_277 TSMC_278 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ S5LLSVTSW8U80_WLDRV4X1 
XMIO_L0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 BWEB[0] BWEB[1] D[0] D[1] Q[0] Q[1] 
+ TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L1 TSMC_13 TSMC_14 TSMC_15 TSMC_16 BWEB[2] BWEB[3] D[2] D[3] Q[2] Q[3] 
+ TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L2 TSMC_17 TSMC_18 TSMC_19 TSMC_20 BWEB[4] BWEB[5] D[4] D[5] Q[4] Q[5] 
+ TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L3 TSMC_21 TSMC_22 TSMC_23 TSMC_24 BWEB[6] BWEB[7] D[6] D[7] Q[6] Q[7] 
+ TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L4 TSMC_25 TSMC_26 TSMC_27 TSMC_28 BWEB[8] BWEB[9] D[8] D[9] Q[8] Q[9] 
+ TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L5 TSMC_29 TSMC_30 TSMC_31 TSMC_32 BWEB[10] BWEB[11] D[10] D[11] Q[10] 
+ Q[11] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L6 TSMC_33 TSMC_34 TSMC_35 TSMC_36 BWEB[12] BWEB[13] D[12] D[13] Q[12] 
+ Q[13] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L7 TSMC_37 TSMC_38 TSMC_39 TSMC_40 BWEB[14] BWEB[15] D[14] D[15] Q[14] 
+ Q[15] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L8 TSMC_41 TSMC_42 TSMC_43 TSMC_44 BWEB[16] BWEB[17] D[16] D[17] Q[16] 
+ Q[17] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L9 TSMC_45 TSMC_46 TSMC_47 TSMC_48 BWEB[18] BWEB[19] D[18] D[19] Q[18] 
+ Q[19] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L10 TSMC_49 TSMC_50 TSMC_51 TSMC_52 BWEB[20] BWEB[21] D[20] D[21] Q[20] 
+ Q[21] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L11 TSMC_53 TSMC_54 TSMC_55 TSMC_56 BWEB[22] BWEB[23] D[22] D[23] Q[22] 
+ Q[23] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L12 TSMC_57 TSMC_58 TSMC_59 TSMC_60 BWEB[24] BWEB[25] D[24] D[25] Q[24] 
+ Q[25] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L13 TSMC_61 TSMC_62 TSMC_63 TSMC_64 BWEB[26] BWEB[27] D[26] D[27] Q[26] 
+ Q[27] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L14 TSMC_65 TSMC_66 TSMC_67 TSMC_68 BWEB[28] BWEB[29] D[28] D[29] Q[28] 
+ Q[29] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L15 TSMC_69 TSMC_70 TSMC_71 TSMC_72 BWEB[30] BWEB[31] D[30] D[31] Q[30] 
+ Q[31] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L16 TSMC_73 TSMC_74 TSMC_75 TSMC_76 BWEB[32] BWEB[33] D[32] D[33] Q[32] 
+ Q[33] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L17 TSMC_77 TSMC_78 TSMC_79 TSMC_80 BWEB[34] BWEB[35] D[34] D[35] Q[34] 
+ Q[35] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L18 TSMC_81 TSMC_82 TSMC_83 TSMC_84 BWEB[36] BWEB[37] D[36] D[37] Q[36] 
+ Q[37] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L19 TSMC_85 TSMC_86 TSMC_87 TSMC_88 BWEB[38] BWEB[39] D[38] D[39] Q[38] 
+ Q[39] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L20 TSMC_89 TSMC_90 TSMC_91 TSMC_92 BWEB[40] BWEB[41] D[40] D[41] Q[40] 
+ Q[41] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L21 TSMC_93 TSMC_94 TSMC_95 TSMC_96 BWEB[42] BWEB[43] D[42] D[43] Q[42] 
+ Q[43] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L22 TSMC_97 TSMC_98 TSMC_99 TSMC_100 BWEB[44] BWEB[45] D[44] D[45] Q[44] 
+ Q[45] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L23 TSMC_101 TSMC_102 TSMC_103 TSMC_104 BWEB[46] BWEB[47] D[46] D[47] 
+ Q[46] Q[47] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L24 TSMC_105 TSMC_106 TSMC_107 TSMC_108 BWEB[48] BWEB[49] D[48] D[49] 
+ Q[48] Q[49] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L25 TSMC_109 TSMC_110 TSMC_111 TSMC_112 BWEB[50] BWEB[51] D[50] D[51] 
+ Q[50] Q[51] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L26 TSMC_113 TSMC_114 TSMC_115 TSMC_116 BWEB[52] BWEB[53] D[52] D[53] 
+ Q[52] Q[53] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L27 TSMC_117 TSMC_118 TSMC_119 TSMC_120 BWEB[54] BWEB[55] D[54] D[55] 
+ Q[54] Q[55] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L28 TSMC_121 TSMC_122 TSMC_123 TSMC_124 BWEB[56] BWEB[57] D[56] D[57] 
+ Q[56] Q[57] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L29 TSMC_125 TSMC_126 TSMC_127 TSMC_128 BWEB[58] BWEB[59] D[58] D[59] 
+ Q[58] Q[59] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L30 TSMC_129 TSMC_130 TSMC_131 TSMC_132 BWEB[60] BWEB[61] D[60] D[61] 
+ Q[60] Q[61] TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_L31 TSMC_133 TSMC_134 TSMC_135 TSMC_136 BWEB[62] BWEB[63] D[62] D[63] 
+ Q[62] Q[63] TSMC_283 TSMC_288 TSMC_289 TSMC_286 TSMC_290 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XIOEDGE_L TSMC_289 TSMC_285 TSMC_286 VDD VDD VSS 
+ S5LLSVTSW8U80_IOEDGE_L_MUX1 
XMIO_R0 TSMC_137 TSMC_138 TSMC_139 TSMC_140 BWEB[64] BWEB[65] D[64] D[65] Q[64] 
+ Q[65] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R1 TSMC_149 TSMC_150 TSMC_151 TSMC_152 BWEB[66] BWEB[67] D[66] D[67] Q[66] 
+ Q[67] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R2 TSMC_153 TSMC_154 TSMC_155 TSMC_156 BWEB[68] BWEB[69] D[68] D[69] Q[68] 
+ Q[69] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R3 TSMC_157 TSMC_158 TSMC_159 TSMC_160 BWEB[70] BWEB[71] D[70] D[71] Q[70] 
+ Q[71] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R4 TSMC_161 TSMC_162 TSMC_163 TSMC_164 BWEB[72] BWEB[73] D[72] D[73] Q[72] 
+ Q[73] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R5 TSMC_165 TSMC_166 TSMC_167 TSMC_168 BWEB[74] BWEB[75] D[74] D[75] Q[74] 
+ Q[75] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R6 TSMC_169 TSMC_170 TSMC_171 TSMC_172 BWEB[76] BWEB[77] D[76] D[77] Q[76] 
+ Q[77] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R7 TSMC_173 TSMC_174 TSMC_175 TSMC_176 BWEB[78] BWEB[79] D[78] D[79] Q[78] 
+ Q[79] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R8 TSMC_177 TSMC_178 TSMC_179 TSMC_180 BWEB[80] BWEB[81] D[80] D[81] Q[80] 
+ Q[81] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R9 TSMC_181 TSMC_182 TSMC_183 TSMC_184 BWEB[82] BWEB[83] D[82] D[83] Q[82] 
+ Q[83] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R10 TSMC_185 TSMC_186 TSMC_187 TSMC_188 BWEB[84] BWEB[85] D[84] D[85] 
+ Q[84] Q[85] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R11 TSMC_189 TSMC_190 TSMC_191 TSMC_192 BWEB[86] BWEB[87] D[86] D[87] 
+ Q[86] Q[87] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R12 TSMC_193 TSMC_194 TSMC_195 TSMC_196 BWEB[88] BWEB[89] D[88] D[89] 
+ Q[88] Q[89] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R13 TSMC_197 TSMC_198 TSMC_199 TSMC_200 BWEB[90] BWEB[91] D[90] D[91] 
+ Q[90] Q[91] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R14 TSMC_201 TSMC_202 TSMC_203 TSMC_204 BWEB[92] BWEB[93] D[92] D[93] 
+ Q[92] Q[93] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R15 TSMC_205 TSMC_206 TSMC_207 TSMC_208 BWEB[94] BWEB[95] D[94] D[95] 
+ Q[94] Q[95] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R16 TSMC_209 TSMC_210 TSMC_211 TSMC_212 BWEB[96] BWEB[97] D[96] D[97] 
+ Q[96] Q[97] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R17 TSMC_213 TSMC_214 TSMC_215 TSMC_216 BWEB[98] BWEB[99] D[98] D[99] 
+ Q[98] Q[99] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R18 TSMC_217 TSMC_218 TSMC_219 TSMC_220 BWEB[100] BWEB[101] D[100] 
+ D[101] Q[100] Q[101] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R19 TSMC_221 TSMC_222 TSMC_223 TSMC_224 BWEB[102] BWEB[103] D[102] 
+ D[103] Q[102] Q[103] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R20 TSMC_225 TSMC_226 TSMC_227 TSMC_228 BWEB[104] BWEB[105] D[104] 
+ D[105] Q[104] Q[105] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R21 TSMC_229 TSMC_230 TSMC_231 TSMC_232 BWEB[106] BWEB[107] D[106] 
+ D[107] Q[106] Q[107] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R22 TSMC_233 TSMC_234 TSMC_235 TSMC_236 BWEB[108] BWEB[109] D[108] 
+ D[109] Q[108] Q[109] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R23 TSMC_237 TSMC_238 TSMC_239 TSMC_240 BWEB[110] BWEB[111] D[110] 
+ D[111] Q[110] Q[111] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R24 TSMC_241 TSMC_242 TSMC_243 TSMC_244 BWEB[112] BWEB[113] D[112] 
+ D[113] Q[112] Q[113] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R25 TSMC_245 TSMC_246 TSMC_247 TSMC_248 BWEB[114] BWEB[115] D[114] 
+ D[115] Q[114] Q[115] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R26 TSMC_249 TSMC_250 TSMC_251 TSMC_252 BWEB[116] BWEB[117] D[116] 
+ D[117] Q[116] Q[117] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R27 TSMC_253 TSMC_254 TSMC_255 TSMC_256 BWEB[118] BWEB[119] D[118] 
+ D[119] Q[118] Q[119] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R28 TSMC_257 TSMC_258 TSMC_259 TSMC_260 BWEB[120] BWEB[121] D[120] 
+ D[121] Q[120] Q[121] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R29 TSMC_261 TSMC_262 TSMC_263 TSMC_264 BWEB[122] BWEB[123] D[122] 
+ D[123] Q[122] Q[123] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R30 TSMC_265 TSMC_266 TSMC_267 TSMC_268 BWEB[124] BWEB[125] D[124] 
+ D[125] Q[124] Q[125] TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XMIO_R31 TSMC_269 TSMC_270 TSMC_271 TSMC_272 BWEB[126] BWEB[127] D[126] 
+ D[127] Q[126] Q[127] TSMC_291 TSMC_296 TSMC_297 TSMC_294 TSMC_298 VDD VSS 
+ S5LLSVTSW8U80_MIO 
XIOEDGE_R TSMC_294 VDD VDD VSS S5LLSVTSW8U80_IOEDGE_R 
XTKBL_CELL_L TSMC_299 TSMC_300 VDD VDD VSS TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 S5LLSVTSW8U80_TKBL_ARR 
XCNT A[0] A[1] A[2] TSMC_301 TSMC_301 TSMC_301 TSMC_301 TSMC_301 CEB TSMC_302 
+ CLK TSMC_301 TSMC_301 TSMC_303 TSMC_304 TSMC_301 TSMC_305 TSMC_306 
+ TSMC_307 TSMC_283 TSMC_291 TSMC_288 TSMC_284 TSMC_292 TSMC_296 
+ TSMC_301 TSMC_308 TSMC_301 TSMC_301 TSMC_301 TSMC_309 TSMC_310 
+ TSMC_311 TSMC_301 TSMC_301 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ TSMC_294 RTSEL[0] RTSEL[1] TSMC_289 TSMC_285 TSMC_293 TSMC_297 
+ TSMC_286 TSMC_301 TSMC_316 TSMC_290 TSMC_287 TSMC_295 TSMC_298 
+ TSMC_301 TSMC_317 TSMC_304 TSMC_301 TSMC_299 TSMC_318 TSMC_300 TSMC_301 VDD 
+ VDD VSS TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_279 TSMC_280 
+ TSMC_281 TSMC_282 TSMC_277 TSMC_319 TSMC_320 TSMC_321 TSMC_278 
+ TSMC_322 TSMC_323 TSMC_324 WEB TSMC_325 TSMC_326 WTSEL[0] WTSEL[1] 
+ S5LLSVTSW8U80_CNTS1_SLP 
XDIOA_A0 A[0] TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_A1 A[1] TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_A2 A[2] TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOBIT_D0 D[0] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_0 BWEB[0] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D1 D[1] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_1 BWEB[1] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D2 D[2] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_2 BWEB[2] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D3 D[3] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_3 BWEB[3] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D4 D[4] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_4 BWEB[4] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D5 D[5] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_5 BWEB[5] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D6 D[6] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_6 BWEB[6] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D7 D[7] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_7 BWEB[7] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D8 D[8] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_8 BWEB[8] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D9 D[9] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_9 BWEB[9] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D10 D[10] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_10 BWEB[10] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D11 D[11] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_11 BWEB[11] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D12 D[12] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_12 BWEB[12] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D13 D[13] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_13 BWEB[13] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D14 D[14] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_14 BWEB[14] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D15 D[15] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_15 BWEB[15] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D16 D[16] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_16 BWEB[16] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D17 D[17] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_17 BWEB[17] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D18 D[18] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_18 BWEB[18] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D19 D[19] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_19 BWEB[19] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D20 D[20] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_20 BWEB[20] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D21 D[21] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_21 BWEB[21] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D22 D[22] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_22 BWEB[22] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D23 D[23] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_23 BWEB[23] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D24 D[24] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_24 BWEB[24] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D25 D[25] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_25 BWEB[25] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D26 D[26] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_26 BWEB[26] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D27 D[27] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_27 BWEB[27] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D28 D[28] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_28 BWEB[28] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D29 D[29] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_29 BWEB[29] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D30 D[30] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_30 BWEB[30] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D31 D[31] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_31 BWEB[31] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D32 D[32] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_32 BWEB[32] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D33 D[33] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_33 BWEB[33] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D34 D[34] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_34 BWEB[34] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D35 D[35] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_35 BWEB[35] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D36 D[36] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_36 BWEB[36] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D37 D[37] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_37 BWEB[37] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D38 D[38] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_38 BWEB[38] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D39 D[39] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_39 BWEB[39] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D40 D[40] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_40 BWEB[40] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D41 D[41] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_41 BWEB[41] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D42 D[42] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_42 BWEB[42] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D43 D[43] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_43 BWEB[43] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D44 D[44] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_44 BWEB[44] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D45 D[45] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_45 BWEB[45] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D46 D[46] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_46 BWEB[46] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D47 D[47] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_47 BWEB[47] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D48 D[48] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_48 BWEB[48] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D49 D[49] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_49 BWEB[49] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D50 D[50] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_50 BWEB[50] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D51 D[51] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_51 BWEB[51] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D52 D[52] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_52 BWEB[52] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D53 D[53] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_53 BWEB[53] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D54 D[54] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_54 BWEB[54] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D55 D[55] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_55 BWEB[55] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D56 D[56] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_56 BWEB[56] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D57 D[57] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_57 BWEB[57] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D58 D[58] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_58 BWEB[58] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D59 D[59] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_59 BWEB[59] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D60 D[60] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_60 BWEB[60] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D61 D[61] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_61 BWEB[61] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D62 D[62] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_62 BWEB[62] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D63 D[63] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_63 BWEB[63] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D64 D[64] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_64 BWEB[64] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D65 D[65] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_65 BWEB[65] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D66 D[66] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_66 BWEB[66] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D67 D[67] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_67 BWEB[67] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D68 D[68] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_68 BWEB[68] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D69 D[69] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_69 BWEB[69] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D70 D[70] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_70 BWEB[70] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D71 D[71] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_71 BWEB[71] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D72 D[72] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_72 BWEB[72] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D73 D[73] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_73 BWEB[73] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D74 D[74] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_74 BWEB[74] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D75 D[75] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_75 BWEB[75] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D76 D[76] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_76 BWEB[76] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D77 D[77] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_77 BWEB[77] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D78 D[78] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_78 BWEB[78] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D79 D[79] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_79 BWEB[79] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D80 D[80] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_80 BWEB[80] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D81 D[81] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_81 BWEB[81] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D82 D[82] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_82 BWEB[82] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D83 D[83] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_83 BWEB[83] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D84 D[84] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_84 BWEB[84] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D85 D[85] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_85 BWEB[85] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D86 D[86] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_86 BWEB[86] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D87 D[87] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_87 BWEB[87] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D88 D[88] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_88 BWEB[88] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D89 D[89] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_89 BWEB[89] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D90 D[90] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_90 BWEB[90] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D91 D[91] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_91 BWEB[91] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D92 D[92] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_92 BWEB[92] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D93 D[93] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_93 BWEB[93] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D94 D[94] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_94 BWEB[94] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D95 D[95] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_95 BWEB[95] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D96 D[96] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_96 BWEB[96] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D97 D[97] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_97 BWEB[97] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D98 D[98] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_98 BWEB[98] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D99 D[99] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_99 BWEB[99] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D100 D[100] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_100 BWEB[100] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D101 D[101] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_101 BWEB[101] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D102 D[102] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_102 BWEB[102] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D103 D[103] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_103 BWEB[103] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D104 D[104] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_104 BWEB[104] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D105 D[105] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_105 BWEB[105] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D106 D[106] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_106 BWEB[106] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D107 D[107] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_107 BWEB[107] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D108 D[108] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_108 BWEB[108] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D109 D[109] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_109 BWEB[109] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D110 D[110] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_110 BWEB[110] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D111 D[111] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_111 BWEB[111] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D112 D[112] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_112 BWEB[112] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D113 D[113] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_113 BWEB[113] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D114 D[114] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_114 BWEB[114] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D115 D[115] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_115 BWEB[115] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D116 D[116] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_116 BWEB[116] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D117 D[117] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_117 BWEB[117] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D118 D[118] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_118 BWEB[118] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D119 D[119] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_119 BWEB[119] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D120 D[120] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_120 BWEB[120] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D121 D[121] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_121 BWEB[121] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D122 D[122] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_122 BWEB[122] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D123 D[123] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_123 BWEB[123] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D124 D[124] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_124 BWEB[124] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D125 D[125] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_125 BWEB[125] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D126 D[126] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_126 BWEB[126] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_D127 D[127] VSS S5LLSVTSW8U80_DIOBIT 
XDIOBIT_BWEB1_127 BWEB[127] VSS S5LLSVTSW8U80_DIOBIT 
XDIOA_WTSEL_0 WTSEL[0] TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_WTSEL_1 WTSEL[1] TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_RTSEL_0 RTSEL[0] TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_RTSEL_1 RTSEL[1] TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_CEB CEB TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_CLK CLK TSMC_301 VSS S5LLSVTSW8U80_DIOA 
XDIOA_WEB WEB TSMC_301 VSS S5LLSVTSW8U80_DIOA 
.ENDS


