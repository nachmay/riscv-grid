# Created by MC2 : Version 2013.12.00.f on 2025/06/23, 08:34:14

#*********************************************************************************************************************/
# Technology     : TSMC 16nm CMOS Logic FinFet Compact (FFC) Low Leakage HKMG                          */
# Memory Type    : TSMC 16nm FFC Single Port SRAM with d0907 bit cell                     */
# Library Name   : ts1n16ffcllsvta64x128m4sw (user specify : ts1n16ffcllsvta64x128m4sw)            */
# Library Version: 120a                                                */
# Generated Time : 2025/06/23, 08:34:08                                        */
#*********************************************************************************************************************/
#                                                            */
# STATEMENT OF USE                                                    */
#                                                            */
# This information contains confidential and proprietary information of TSMC.                    */
# No part of this information may be reproduced, transmitted, transcribed,                        */
# stored in a retrieval system, or translated into any human or computer                        */
# language, in any form or by any means, electronic, mechanical, magnetic,                        */
# optical, chemical, manual, or otherwise, without the prior written permission                    */
# of TSMC. This information was prepared for informational purpose and is for                    */
# use by TSMC's customers only. TSMC reserves the right to make changes in the                    */
# information at any time and without notice.                                    */
#                                                            */
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N16FFCLLSVTA64X128M4SW
	CLASS BLOCK ;
	FOREIGN TS1N16FFCLLSVTA64X128M4SW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 17.375 BY 272.880 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 131.720 17.375 131.800 ;
			LAYER M2 ;
			RECT 17.127 131.720 17.375 131.800 ;
			LAYER M3 ;
			RECT 17.127 131.720 17.375 131.800 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 130.376 17.375 130.456 ;
			LAYER M2 ;
			RECT 17.127 130.376 17.375 130.456 ;
			LAYER M3 ;
			RECT 17.127 130.376 17.375 130.456 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 140.744 17.375 140.824 ;
			LAYER M2 ;
			RECT 17.127 140.744 17.375 140.824 ;
			LAYER M3 ;
			RECT 17.127 140.744 17.375 140.824 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 139.976 17.375 140.056 ;
			LAYER M2 ;
			RECT 17.127 139.976 17.375 140.056 ;
			LAYER M3 ;
			RECT 17.127 139.976 17.375 140.056 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 139.400 17.375 139.480 ;
			LAYER M2 ;
			RECT 17.127 139.400 17.375 139.480 ;
			LAYER M3 ;
			RECT 17.127 139.400 17.375 139.480 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 136.712 17.375 136.792 ;
			LAYER M2 ;
			RECT 17.127 136.712 17.375 136.792 ;
			LAYER M3 ;
			RECT 17.127 136.712 17.375 136.792 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[5]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 1.976 17.375 2.056 ;
			LAYER M2 ;
			RECT 17.127 1.976 17.375 2.056 ;
			LAYER M3 ;
			RECT 17.127 1.976 17.375 2.056 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 3.992 17.375 4.072 ;
			LAYER M2 ;
			RECT 17.127 3.992 17.375 4.072 ;
			LAYER M3 ;
			RECT 17.127 3.992 17.375 4.072 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 6.008 17.375 6.088 ;
			LAYER M2 ;
			RECT 17.127 6.008 17.375 6.088 ;
			LAYER M3 ;
			RECT 17.127 6.008 17.375 6.088 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 8.024 17.375 8.104 ;
			LAYER M2 ;
			RECT 17.127 8.024 17.375 8.104 ;
			LAYER M3 ;
			RECT 17.127 8.024 17.375 8.104 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 10.040 17.375 10.120 ;
			LAYER M2 ;
			RECT 17.127 10.040 17.375 10.120 ;
			LAYER M3 ;
			RECT 17.127 10.040 17.375 10.120 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 12.056 17.375 12.136 ;
			LAYER M2 ;
			RECT 17.127 12.056 17.375 12.136 ;
			LAYER M3 ;
			RECT 17.127 12.056 17.375 12.136 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 14.072 17.375 14.152 ;
			LAYER M2 ;
			RECT 17.127 14.072 17.375 14.152 ;
			LAYER M3 ;
			RECT 17.127 14.072 17.375 14.152 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 16.088 17.375 16.168 ;
			LAYER M2 ;
			RECT 17.127 16.088 17.375 16.168 ;
			LAYER M3 ;
			RECT 17.127 16.088 17.375 16.168 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 18.104 17.375 18.184 ;
			LAYER M2 ;
			RECT 17.127 18.104 17.375 18.184 ;
			LAYER M3 ;
			RECT 17.127 18.104 17.375 18.184 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 20.120 17.375 20.200 ;
			LAYER M2 ;
			RECT 17.127 20.120 17.375 20.200 ;
			LAYER M3 ;
			RECT 17.127 20.120 17.375 20.200 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 22.136 17.375 22.216 ;
			LAYER M2 ;
			RECT 17.127 22.136 17.375 22.216 ;
			LAYER M3 ;
			RECT 17.127 22.136 17.375 22.216 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 24.152 17.375 24.232 ;
			LAYER M2 ;
			RECT 17.127 24.152 17.375 24.232 ;
			LAYER M3 ;
			RECT 17.127 24.152 17.375 24.232 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 26.168 17.375 26.248 ;
			LAYER M2 ;
			RECT 17.127 26.168 17.375 26.248 ;
			LAYER M3 ;
			RECT 17.127 26.168 17.375 26.248 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 28.184 17.375 28.264 ;
			LAYER M2 ;
			RECT 17.127 28.184 17.375 28.264 ;
			LAYER M3 ;
			RECT 17.127 28.184 17.375 28.264 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 30.200 17.375 30.280 ;
			LAYER M2 ;
			RECT 17.127 30.200 17.375 30.280 ;
			LAYER M3 ;
			RECT 17.127 30.200 17.375 30.280 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 32.216 17.375 32.296 ;
			LAYER M2 ;
			RECT 17.127 32.216 17.375 32.296 ;
			LAYER M3 ;
			RECT 17.127 32.216 17.375 32.296 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 34.232 17.375 34.312 ;
			LAYER M2 ;
			RECT 17.127 34.232 17.375 34.312 ;
			LAYER M3 ;
			RECT 17.127 34.232 17.375 34.312 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 36.248 17.375 36.328 ;
			LAYER M2 ;
			RECT 17.127 36.248 17.375 36.328 ;
			LAYER M3 ;
			RECT 17.127 36.248 17.375 36.328 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 38.264 17.375 38.344 ;
			LAYER M2 ;
			RECT 17.127 38.264 17.375 38.344 ;
			LAYER M3 ;
			RECT 17.127 38.264 17.375 38.344 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 40.280 17.375 40.360 ;
			LAYER M2 ;
			RECT 17.127 40.280 17.375 40.360 ;
			LAYER M3 ;
			RECT 17.127 40.280 17.375 40.360 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 42.296 17.375 42.376 ;
			LAYER M2 ;
			RECT 17.127 42.296 17.375 42.376 ;
			LAYER M3 ;
			RECT 17.127 42.296 17.375 42.376 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 44.312 17.375 44.392 ;
			LAYER M2 ;
			RECT 17.127 44.312 17.375 44.392 ;
			LAYER M3 ;
			RECT 17.127 44.312 17.375 44.392 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 46.328 17.375 46.408 ;
			LAYER M2 ;
			RECT 17.127 46.328 17.375 46.408 ;
			LAYER M3 ;
			RECT 17.127 46.328 17.375 46.408 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 48.344 17.375 48.424 ;
			LAYER M2 ;
			RECT 17.127 48.344 17.375 48.424 ;
			LAYER M3 ;
			RECT 17.127 48.344 17.375 48.424 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 50.360 17.375 50.440 ;
			LAYER M2 ;
			RECT 17.127 50.360 17.375 50.440 ;
			LAYER M3 ;
			RECT 17.127 50.360 17.375 50.440 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 52.376 17.375 52.456 ;
			LAYER M2 ;
			RECT 17.127 52.376 17.375 52.456 ;
			LAYER M3 ;
			RECT 17.127 52.376 17.375 52.456 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 54.392 17.375 54.472 ;
			LAYER M2 ;
			RECT 17.127 54.392 17.375 54.472 ;
			LAYER M3 ;
			RECT 17.127 54.392 17.375 54.472 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 56.408 17.375 56.488 ;
			LAYER M2 ;
			RECT 17.127 56.408 17.375 56.488 ;
			LAYER M3 ;
			RECT 17.127 56.408 17.375 56.488 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 58.424 17.375 58.504 ;
			LAYER M2 ;
			RECT 17.127 58.424 17.375 58.504 ;
			LAYER M3 ;
			RECT 17.127 58.424 17.375 58.504 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 60.440 17.375 60.520 ;
			LAYER M2 ;
			RECT 17.127 60.440 17.375 60.520 ;
			LAYER M3 ;
			RECT 17.127 60.440 17.375 60.520 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 62.456 17.375 62.536 ;
			LAYER M2 ;
			RECT 17.127 62.456 17.375 62.536 ;
			LAYER M3 ;
			RECT 17.127 62.456 17.375 62.536 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 64.472 17.375 64.552 ;
			LAYER M2 ;
			RECT 17.127 64.472 17.375 64.552 ;
			LAYER M3 ;
			RECT 17.127 64.472 17.375 64.552 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[31]

	PIN BWEB[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 66.488 17.375 66.568 ;
			LAYER M2 ;
			RECT 17.127 66.488 17.375 66.568 ;
			LAYER M3 ;
			RECT 17.127 66.488 17.375 66.568 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[32]

	PIN BWEB[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 68.504 17.375 68.584 ;
			LAYER M2 ;
			RECT 17.127 68.504 17.375 68.584 ;
			LAYER M3 ;
			RECT 17.127 68.504 17.375 68.584 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[33]

	PIN BWEB[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 70.520 17.375 70.600 ;
			LAYER M2 ;
			RECT 17.127 70.520 17.375 70.600 ;
			LAYER M3 ;
			RECT 17.127 70.520 17.375 70.600 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[34]

	PIN BWEB[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 72.536 17.375 72.616 ;
			LAYER M2 ;
			RECT 17.127 72.536 17.375 72.616 ;
			LAYER M3 ;
			RECT 17.127 72.536 17.375 72.616 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[35]

	PIN BWEB[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 74.552 17.375 74.632 ;
			LAYER M2 ;
			RECT 17.127 74.552 17.375 74.632 ;
			LAYER M3 ;
			RECT 17.127 74.552 17.375 74.632 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[36]

	PIN BWEB[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 76.568 17.375 76.648 ;
			LAYER M2 ;
			RECT 17.127 76.568 17.375 76.648 ;
			LAYER M3 ;
			RECT 17.127 76.568 17.375 76.648 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[37]

	PIN BWEB[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 78.584 17.375 78.664 ;
			LAYER M2 ;
			RECT 17.127 78.584 17.375 78.664 ;
			LAYER M3 ;
			RECT 17.127 78.584 17.375 78.664 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[38]

	PIN BWEB[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 80.600 17.375 80.680 ;
			LAYER M2 ;
			RECT 17.127 80.600 17.375 80.680 ;
			LAYER M3 ;
			RECT 17.127 80.600 17.375 80.680 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[39]

	PIN BWEB[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 82.616 17.375 82.696 ;
			LAYER M2 ;
			RECT 17.127 82.616 17.375 82.696 ;
			LAYER M3 ;
			RECT 17.127 82.616 17.375 82.696 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[40]

	PIN BWEB[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 84.632 17.375 84.712 ;
			LAYER M2 ;
			RECT 17.127 84.632 17.375 84.712 ;
			LAYER M3 ;
			RECT 17.127 84.632 17.375 84.712 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[41]

	PIN BWEB[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 86.648 17.375 86.728 ;
			LAYER M2 ;
			RECT 17.127 86.648 17.375 86.728 ;
			LAYER M3 ;
			RECT 17.127 86.648 17.375 86.728 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[42]

	PIN BWEB[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 88.664 17.375 88.744 ;
			LAYER M2 ;
			RECT 17.127 88.664 17.375 88.744 ;
			LAYER M3 ;
			RECT 17.127 88.664 17.375 88.744 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[43]

	PIN BWEB[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 90.680 17.375 90.760 ;
			LAYER M2 ;
			RECT 17.127 90.680 17.375 90.760 ;
			LAYER M3 ;
			RECT 17.127 90.680 17.375 90.760 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[44]

	PIN BWEB[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 92.696 17.375 92.776 ;
			LAYER M2 ;
			RECT 17.127 92.696 17.375 92.776 ;
			LAYER M3 ;
			RECT 17.127 92.696 17.375 92.776 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[45]

	PIN BWEB[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 94.712 17.375 94.792 ;
			LAYER M2 ;
			RECT 17.127 94.712 17.375 94.792 ;
			LAYER M3 ;
			RECT 17.127 94.712 17.375 94.792 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[46]

	PIN BWEB[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 96.728 17.375 96.808 ;
			LAYER M2 ;
			RECT 17.127 96.728 17.375 96.808 ;
			LAYER M3 ;
			RECT 17.127 96.728 17.375 96.808 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[47]

	PIN BWEB[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 98.744 17.375 98.824 ;
			LAYER M2 ;
			RECT 17.127 98.744 17.375 98.824 ;
			LAYER M3 ;
			RECT 17.127 98.744 17.375 98.824 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[48]

	PIN BWEB[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 100.760 17.375 100.840 ;
			LAYER M2 ;
			RECT 17.127 100.760 17.375 100.840 ;
			LAYER M3 ;
			RECT 17.127 100.760 17.375 100.840 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[49]

	PIN BWEB[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 102.776 17.375 102.856 ;
			LAYER M2 ;
			RECT 17.127 102.776 17.375 102.856 ;
			LAYER M3 ;
			RECT 17.127 102.776 17.375 102.856 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[50]

	PIN BWEB[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 104.792 17.375 104.872 ;
			LAYER M2 ;
			RECT 17.127 104.792 17.375 104.872 ;
			LAYER M3 ;
			RECT 17.127 104.792 17.375 104.872 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[51]

	PIN BWEB[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 106.808 17.375 106.888 ;
			LAYER M2 ;
			RECT 17.127 106.808 17.375 106.888 ;
			LAYER M3 ;
			RECT 17.127 106.808 17.375 106.888 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[52]

	PIN BWEB[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 108.824 17.375 108.904 ;
			LAYER M2 ;
			RECT 17.127 108.824 17.375 108.904 ;
			LAYER M3 ;
			RECT 17.127 108.824 17.375 108.904 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[53]

	PIN BWEB[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 110.840 17.375 110.920 ;
			LAYER M2 ;
			RECT 17.127 110.840 17.375 110.920 ;
			LAYER M3 ;
			RECT 17.127 110.840 17.375 110.920 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[54]

	PIN BWEB[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 112.856 17.375 112.936 ;
			LAYER M2 ;
			RECT 17.127 112.856 17.375 112.936 ;
			LAYER M3 ;
			RECT 17.127 112.856 17.375 112.936 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[55]

	PIN BWEB[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 114.872 17.375 114.952 ;
			LAYER M2 ;
			RECT 17.127 114.872 17.375 114.952 ;
			LAYER M3 ;
			RECT 17.127 114.872 17.375 114.952 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[56]

	PIN BWEB[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 116.888 17.375 116.968 ;
			LAYER M2 ;
			RECT 17.127 116.888 17.375 116.968 ;
			LAYER M3 ;
			RECT 17.127 116.888 17.375 116.968 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[57]

	PIN BWEB[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 118.904 17.375 118.984 ;
			LAYER M2 ;
			RECT 17.127 118.904 17.375 118.984 ;
			LAYER M3 ;
			RECT 17.127 118.904 17.375 118.984 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[58]

	PIN BWEB[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 120.920 17.375 121.000 ;
			LAYER M2 ;
			RECT 17.127 120.920 17.375 121.000 ;
			LAYER M3 ;
			RECT 17.127 120.920 17.375 121.000 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[59]

	PIN BWEB[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 122.936 17.375 123.016 ;
			LAYER M2 ;
			RECT 17.127 122.936 17.375 123.016 ;
			LAYER M3 ;
			RECT 17.127 122.936 17.375 123.016 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[60]

	PIN BWEB[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 124.952 17.375 125.032 ;
			LAYER M2 ;
			RECT 17.127 124.952 17.375 125.032 ;
			LAYER M3 ;
			RECT 17.127 124.952 17.375 125.032 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[61]

	PIN BWEB[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 126.968 17.375 127.048 ;
			LAYER M2 ;
			RECT 17.127 126.968 17.375 127.048 ;
			LAYER M3 ;
			RECT 17.127 126.968 17.375 127.048 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[62]

	PIN BWEB[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 128.984 17.375 129.064 ;
			LAYER M2 ;
			RECT 17.127 128.984 17.375 129.064 ;
			LAYER M3 ;
			RECT 17.127 128.984 17.375 129.064 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[63]

	PIN BWEB[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 143.864 17.375 143.944 ;
			LAYER M2 ;
			RECT 17.127 143.864 17.375 143.944 ;
			LAYER M3 ;
			RECT 17.127 143.864 17.375 143.944 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[64]

	PIN BWEB[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 145.880 17.375 145.960 ;
			LAYER M2 ;
			RECT 17.127 145.880 17.375 145.960 ;
			LAYER M3 ;
			RECT 17.127 145.880 17.375 145.960 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[65]

	PIN BWEB[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 147.896 17.375 147.976 ;
			LAYER M2 ;
			RECT 17.127 147.896 17.375 147.976 ;
			LAYER M3 ;
			RECT 17.127 147.896 17.375 147.976 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[66]

	PIN BWEB[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 149.912 17.375 149.992 ;
			LAYER M2 ;
			RECT 17.127 149.912 17.375 149.992 ;
			LAYER M3 ;
			RECT 17.127 149.912 17.375 149.992 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[67]

	PIN BWEB[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 151.928 17.375 152.008 ;
			LAYER M2 ;
			RECT 17.127 151.928 17.375 152.008 ;
			LAYER M3 ;
			RECT 17.127 151.928 17.375 152.008 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[68]

	PIN BWEB[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 153.944 17.375 154.024 ;
			LAYER M2 ;
			RECT 17.127 153.944 17.375 154.024 ;
			LAYER M3 ;
			RECT 17.127 153.944 17.375 154.024 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[69]

	PIN BWEB[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 155.960 17.375 156.040 ;
			LAYER M2 ;
			RECT 17.127 155.960 17.375 156.040 ;
			LAYER M3 ;
			RECT 17.127 155.960 17.375 156.040 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[70]

	PIN BWEB[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 157.976 17.375 158.056 ;
			LAYER M2 ;
			RECT 17.127 157.976 17.375 158.056 ;
			LAYER M3 ;
			RECT 17.127 157.976 17.375 158.056 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[71]

	PIN BWEB[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 159.992 17.375 160.072 ;
			LAYER M2 ;
			RECT 17.127 159.992 17.375 160.072 ;
			LAYER M3 ;
			RECT 17.127 159.992 17.375 160.072 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[72]

	PIN BWEB[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 162.008 17.375 162.088 ;
			LAYER M2 ;
			RECT 17.127 162.008 17.375 162.088 ;
			LAYER M3 ;
			RECT 17.127 162.008 17.375 162.088 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[73]

	PIN BWEB[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 164.024 17.375 164.104 ;
			LAYER M2 ;
			RECT 17.127 164.024 17.375 164.104 ;
			LAYER M3 ;
			RECT 17.127 164.024 17.375 164.104 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[74]

	PIN BWEB[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 166.040 17.375 166.120 ;
			LAYER M2 ;
			RECT 17.127 166.040 17.375 166.120 ;
			LAYER M3 ;
			RECT 17.127 166.040 17.375 166.120 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[75]

	PIN BWEB[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 168.056 17.375 168.136 ;
			LAYER M2 ;
			RECT 17.127 168.056 17.375 168.136 ;
			LAYER M3 ;
			RECT 17.127 168.056 17.375 168.136 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[76]

	PIN BWEB[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 170.072 17.375 170.152 ;
			LAYER M2 ;
			RECT 17.127 170.072 17.375 170.152 ;
			LAYER M3 ;
			RECT 17.127 170.072 17.375 170.152 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[77]

	PIN BWEB[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 172.088 17.375 172.168 ;
			LAYER M2 ;
			RECT 17.127 172.088 17.375 172.168 ;
			LAYER M3 ;
			RECT 17.127 172.088 17.375 172.168 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[78]

	PIN BWEB[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 174.104 17.375 174.184 ;
			LAYER M2 ;
			RECT 17.127 174.104 17.375 174.184 ;
			LAYER M3 ;
			RECT 17.127 174.104 17.375 174.184 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[79]

	PIN BWEB[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 176.120 17.375 176.200 ;
			LAYER M2 ;
			RECT 17.127 176.120 17.375 176.200 ;
			LAYER M3 ;
			RECT 17.127 176.120 17.375 176.200 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[80]

	PIN BWEB[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 178.136 17.375 178.216 ;
			LAYER M2 ;
			RECT 17.127 178.136 17.375 178.216 ;
			LAYER M3 ;
			RECT 17.127 178.136 17.375 178.216 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[81]

	PIN BWEB[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 180.152 17.375 180.232 ;
			LAYER M2 ;
			RECT 17.127 180.152 17.375 180.232 ;
			LAYER M3 ;
			RECT 17.127 180.152 17.375 180.232 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[82]

	PIN BWEB[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 182.168 17.375 182.248 ;
			LAYER M2 ;
			RECT 17.127 182.168 17.375 182.248 ;
			LAYER M3 ;
			RECT 17.127 182.168 17.375 182.248 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[83]

	PIN BWEB[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 184.184 17.375 184.264 ;
			LAYER M2 ;
			RECT 17.127 184.184 17.375 184.264 ;
			LAYER M3 ;
			RECT 17.127 184.184 17.375 184.264 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[84]

	PIN BWEB[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 186.200 17.375 186.280 ;
			LAYER M2 ;
			RECT 17.127 186.200 17.375 186.280 ;
			LAYER M3 ;
			RECT 17.127 186.200 17.375 186.280 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[85]

	PIN BWEB[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 188.216 17.375 188.296 ;
			LAYER M2 ;
			RECT 17.127 188.216 17.375 188.296 ;
			LAYER M3 ;
			RECT 17.127 188.216 17.375 188.296 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[86]

	PIN BWEB[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 190.232 17.375 190.312 ;
			LAYER M2 ;
			RECT 17.127 190.232 17.375 190.312 ;
			LAYER M3 ;
			RECT 17.127 190.232 17.375 190.312 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[87]

	PIN BWEB[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 192.248 17.375 192.328 ;
			LAYER M2 ;
			RECT 17.127 192.248 17.375 192.328 ;
			LAYER M3 ;
			RECT 17.127 192.248 17.375 192.328 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[88]

	PIN BWEB[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 194.264 17.375 194.344 ;
			LAYER M2 ;
			RECT 17.127 194.264 17.375 194.344 ;
			LAYER M3 ;
			RECT 17.127 194.264 17.375 194.344 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[89]

	PIN BWEB[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 196.280 17.375 196.360 ;
			LAYER M2 ;
			RECT 17.127 196.280 17.375 196.360 ;
			LAYER M3 ;
			RECT 17.127 196.280 17.375 196.360 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[90]

	PIN BWEB[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 198.296 17.375 198.376 ;
			LAYER M2 ;
			RECT 17.127 198.296 17.375 198.376 ;
			LAYER M3 ;
			RECT 17.127 198.296 17.375 198.376 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[91]

	PIN BWEB[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 200.312 17.375 200.392 ;
			LAYER M2 ;
			RECT 17.127 200.312 17.375 200.392 ;
			LAYER M3 ;
			RECT 17.127 200.312 17.375 200.392 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[92]

	PIN BWEB[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 202.328 17.375 202.408 ;
			LAYER M2 ;
			RECT 17.127 202.328 17.375 202.408 ;
			LAYER M3 ;
			RECT 17.127 202.328 17.375 202.408 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[93]

	PIN BWEB[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 204.344 17.375 204.424 ;
			LAYER M2 ;
			RECT 17.127 204.344 17.375 204.424 ;
			LAYER M3 ;
			RECT 17.127 204.344 17.375 204.424 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[94]

	PIN BWEB[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 206.360 17.375 206.440 ;
			LAYER M2 ;
			RECT 17.127 206.360 17.375 206.440 ;
			LAYER M3 ;
			RECT 17.127 206.360 17.375 206.440 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[95]

	PIN BWEB[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 208.376 17.375 208.456 ;
			LAYER M2 ;
			RECT 17.127 208.376 17.375 208.456 ;
			LAYER M3 ;
			RECT 17.127 208.376 17.375 208.456 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[96]

	PIN BWEB[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 210.392 17.375 210.472 ;
			LAYER M2 ;
			RECT 17.127 210.392 17.375 210.472 ;
			LAYER M3 ;
			RECT 17.127 210.392 17.375 210.472 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[97]

	PIN BWEB[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 212.408 17.375 212.488 ;
			LAYER M2 ;
			RECT 17.127 212.408 17.375 212.488 ;
			LAYER M3 ;
			RECT 17.127 212.408 17.375 212.488 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[98]

	PIN BWEB[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 214.424 17.375 214.504 ;
			LAYER M2 ;
			RECT 17.127 214.424 17.375 214.504 ;
			LAYER M3 ;
			RECT 17.127 214.424 17.375 214.504 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[99]

	PIN BWEB[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 216.440 17.375 216.520 ;
			LAYER M2 ;
			RECT 17.127 216.440 17.375 216.520 ;
			LAYER M3 ;
			RECT 17.127 216.440 17.375 216.520 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[100]

	PIN BWEB[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 218.456 17.375 218.536 ;
			LAYER M2 ;
			RECT 17.127 218.456 17.375 218.536 ;
			LAYER M3 ;
			RECT 17.127 218.456 17.375 218.536 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[101]

	PIN BWEB[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 220.472 17.375 220.552 ;
			LAYER M2 ;
			RECT 17.127 220.472 17.375 220.552 ;
			LAYER M3 ;
			RECT 17.127 220.472 17.375 220.552 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[102]

	PIN BWEB[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 222.488 17.375 222.568 ;
			LAYER M2 ;
			RECT 17.127 222.488 17.375 222.568 ;
			LAYER M3 ;
			RECT 17.127 222.488 17.375 222.568 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[103]

	PIN BWEB[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 224.504 17.375 224.584 ;
			LAYER M2 ;
			RECT 17.127 224.504 17.375 224.584 ;
			LAYER M3 ;
			RECT 17.127 224.504 17.375 224.584 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[104]

	PIN BWEB[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 226.520 17.375 226.600 ;
			LAYER M2 ;
			RECT 17.127 226.520 17.375 226.600 ;
			LAYER M3 ;
			RECT 17.127 226.520 17.375 226.600 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[105]

	PIN BWEB[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 228.536 17.375 228.616 ;
			LAYER M2 ;
			RECT 17.127 228.536 17.375 228.616 ;
			LAYER M3 ;
			RECT 17.127 228.536 17.375 228.616 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[106]

	PIN BWEB[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 230.552 17.375 230.632 ;
			LAYER M2 ;
			RECT 17.127 230.552 17.375 230.632 ;
			LAYER M3 ;
			RECT 17.127 230.552 17.375 230.632 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[107]

	PIN BWEB[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 232.568 17.375 232.648 ;
			LAYER M2 ;
			RECT 17.127 232.568 17.375 232.648 ;
			LAYER M3 ;
			RECT 17.127 232.568 17.375 232.648 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[108]

	PIN BWEB[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 234.584 17.375 234.664 ;
			LAYER M2 ;
			RECT 17.127 234.584 17.375 234.664 ;
			LAYER M3 ;
			RECT 17.127 234.584 17.375 234.664 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[109]

	PIN BWEB[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 236.600 17.375 236.680 ;
			LAYER M2 ;
			RECT 17.127 236.600 17.375 236.680 ;
			LAYER M3 ;
			RECT 17.127 236.600 17.375 236.680 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[110]

	PIN BWEB[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 238.616 17.375 238.696 ;
			LAYER M2 ;
			RECT 17.127 238.616 17.375 238.696 ;
			LAYER M3 ;
			RECT 17.127 238.616 17.375 238.696 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[111]

	PIN BWEB[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 240.632 17.375 240.712 ;
			LAYER M2 ;
			RECT 17.127 240.632 17.375 240.712 ;
			LAYER M3 ;
			RECT 17.127 240.632 17.375 240.712 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[112]

	PIN BWEB[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 242.648 17.375 242.728 ;
			LAYER M2 ;
			RECT 17.127 242.648 17.375 242.728 ;
			LAYER M3 ;
			RECT 17.127 242.648 17.375 242.728 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[113]

	PIN BWEB[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 244.664 17.375 244.744 ;
			LAYER M2 ;
			RECT 17.127 244.664 17.375 244.744 ;
			LAYER M3 ;
			RECT 17.127 244.664 17.375 244.744 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[114]

	PIN BWEB[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 246.680 17.375 246.760 ;
			LAYER M2 ;
			RECT 17.127 246.680 17.375 246.760 ;
			LAYER M3 ;
			RECT 17.127 246.680 17.375 246.760 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[115]

	PIN BWEB[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 248.696 17.375 248.776 ;
			LAYER M2 ;
			RECT 17.127 248.696 17.375 248.776 ;
			LAYER M3 ;
			RECT 17.127 248.696 17.375 248.776 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[116]

	PIN BWEB[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 250.712 17.375 250.792 ;
			LAYER M2 ;
			RECT 17.127 250.712 17.375 250.792 ;
			LAYER M3 ;
			RECT 17.127 250.712 17.375 250.792 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[117]

	PIN BWEB[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 252.728 17.375 252.808 ;
			LAYER M2 ;
			RECT 17.127 252.728 17.375 252.808 ;
			LAYER M3 ;
			RECT 17.127 252.728 17.375 252.808 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[118]

	PIN BWEB[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 254.744 17.375 254.824 ;
			LAYER M2 ;
			RECT 17.127 254.744 17.375 254.824 ;
			LAYER M3 ;
			RECT 17.127 254.744 17.375 254.824 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[119]

	PIN BWEB[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 256.760 17.375 256.840 ;
			LAYER M2 ;
			RECT 17.127 256.760 17.375 256.840 ;
			LAYER M3 ;
			RECT 17.127 256.760 17.375 256.840 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[120]

	PIN BWEB[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 258.776 17.375 258.856 ;
			LAYER M2 ;
			RECT 17.127 258.776 17.375 258.856 ;
			LAYER M3 ;
			RECT 17.127 258.776 17.375 258.856 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[121]

	PIN BWEB[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 260.792 17.375 260.872 ;
			LAYER M2 ;
			RECT 17.127 260.792 17.375 260.872 ;
			LAYER M3 ;
			RECT 17.127 260.792 17.375 260.872 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[122]

	PIN BWEB[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 262.808 17.375 262.888 ;
			LAYER M2 ;
			RECT 17.127 262.808 17.375 262.888 ;
			LAYER M3 ;
			RECT 17.127 262.808 17.375 262.888 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[123]

	PIN BWEB[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 264.824 17.375 264.904 ;
			LAYER M2 ;
			RECT 17.127 264.824 17.375 264.904 ;
			LAYER M3 ;
			RECT 17.127 264.824 17.375 264.904 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[124]

	PIN BWEB[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 266.840 17.375 266.920 ;
			LAYER M2 ;
			RECT 17.127 266.840 17.375 266.920 ;
			LAYER M3 ;
			RECT 17.127 266.840 17.375 266.920 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[125]

	PIN BWEB[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 268.856 17.375 268.936 ;
			LAYER M2 ;
			RECT 17.127 268.856 17.375 268.936 ;
			LAYER M3 ;
			RECT 17.127 268.856 17.375 268.936 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[126]

	PIN BWEB[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 270.872 17.375 270.952 ;
			LAYER M2 ;
			RECT 17.127 270.872 17.375 270.952 ;
			LAYER M3 ;
			RECT 17.127 270.872 17.375 270.952 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[127]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 133.448 17.375 133.528 ;
			LAYER M2 ;
			RECT 17.127 133.448 17.375 133.528 ;
			LAYER M3 ;
			RECT 17.127 133.448 17.375 133.528 ;
		END
		ANTENNAGATEAREA 0.010000 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081400 LAYER M1 ;
		ANTENNAMAXAREACAR 2.270000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.204800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010000 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.590000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.409600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010000 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.158200 LAYER M3 ;
		ANTENNAMAXAREACAR 25.420000 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 135.752 17.375 135.832 ;
			LAYER M2 ;
			RECT 17.127 135.752 17.375 135.832 ;
			LAYER M3 ;
			RECT 17.127 135.752 17.375 135.832 ;
		END
		ANTENNAGATEAREA 0.284200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 2.071400 LAYER M1 ;
		ANTENNAMAXAREACAR 12.657200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.061400 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.284200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 3.218800 LAYER M2 ;
		ANTENNAMAXAREACAR 73.469000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.031800 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.789800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.284200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.817000 LAYER M3 ;
		ANTENNAMAXAREACAR 83.379800 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 2.360 17.375 2.440 ;
			LAYER M2 ;
			RECT 17.127 2.360 17.375 2.440 ;
			LAYER M3 ;
			RECT 17.127 2.360 17.375 2.440 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 4.376 17.375 4.456 ;
			LAYER M2 ;
			RECT 17.127 4.376 17.375 4.456 ;
			LAYER M3 ;
			RECT 17.127 4.376 17.375 4.456 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 6.392 17.375 6.472 ;
			LAYER M2 ;
			RECT 17.127 6.392 17.375 6.472 ;
			LAYER M3 ;
			RECT 17.127 6.392 17.375 6.472 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 8.408 17.375 8.488 ;
			LAYER M2 ;
			RECT 17.127 8.408 17.375 8.488 ;
			LAYER M3 ;
			RECT 17.127 8.408 17.375 8.488 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 10.424 17.375 10.504 ;
			LAYER M2 ;
			RECT 17.127 10.424 17.375 10.504 ;
			LAYER M3 ;
			RECT 17.127 10.424 17.375 10.504 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 12.440 17.375 12.520 ;
			LAYER M2 ;
			RECT 17.127 12.440 17.375 12.520 ;
			LAYER M3 ;
			RECT 17.127 12.440 17.375 12.520 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 14.456 17.375 14.536 ;
			LAYER M2 ;
			RECT 17.127 14.456 17.375 14.536 ;
			LAYER M3 ;
			RECT 17.127 14.456 17.375 14.536 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 16.472 17.375 16.552 ;
			LAYER M2 ;
			RECT 17.127 16.472 17.375 16.552 ;
			LAYER M3 ;
			RECT 17.127 16.472 17.375 16.552 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 18.488 17.375 18.568 ;
			LAYER M2 ;
			RECT 17.127 18.488 17.375 18.568 ;
			LAYER M3 ;
			RECT 17.127 18.488 17.375 18.568 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 20.504 17.375 20.584 ;
			LAYER M2 ;
			RECT 17.127 20.504 17.375 20.584 ;
			LAYER M3 ;
			RECT 17.127 20.504 17.375 20.584 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 22.520 17.375 22.600 ;
			LAYER M2 ;
			RECT 17.127 22.520 17.375 22.600 ;
			LAYER M3 ;
			RECT 17.127 22.520 17.375 22.600 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 24.536 17.375 24.616 ;
			LAYER M2 ;
			RECT 17.127 24.536 17.375 24.616 ;
			LAYER M3 ;
			RECT 17.127 24.536 17.375 24.616 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 26.552 17.375 26.632 ;
			LAYER M2 ;
			RECT 17.127 26.552 17.375 26.632 ;
			LAYER M3 ;
			RECT 17.127 26.552 17.375 26.632 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 28.568 17.375 28.648 ;
			LAYER M2 ;
			RECT 17.127 28.568 17.375 28.648 ;
			LAYER M3 ;
			RECT 17.127 28.568 17.375 28.648 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 30.584 17.375 30.664 ;
			LAYER M2 ;
			RECT 17.127 30.584 17.375 30.664 ;
			LAYER M3 ;
			RECT 17.127 30.584 17.375 30.664 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 32.600 17.375 32.680 ;
			LAYER M2 ;
			RECT 17.127 32.600 17.375 32.680 ;
			LAYER M3 ;
			RECT 17.127 32.600 17.375 32.680 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 34.616 17.375 34.696 ;
			LAYER M2 ;
			RECT 17.127 34.616 17.375 34.696 ;
			LAYER M3 ;
			RECT 17.127 34.616 17.375 34.696 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 36.632 17.375 36.712 ;
			LAYER M2 ;
			RECT 17.127 36.632 17.375 36.712 ;
			LAYER M3 ;
			RECT 17.127 36.632 17.375 36.712 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 38.648 17.375 38.728 ;
			LAYER M2 ;
			RECT 17.127 38.648 17.375 38.728 ;
			LAYER M3 ;
			RECT 17.127 38.648 17.375 38.728 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 40.664 17.375 40.744 ;
			LAYER M2 ;
			RECT 17.127 40.664 17.375 40.744 ;
			LAYER M3 ;
			RECT 17.127 40.664 17.375 40.744 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 42.680 17.375 42.760 ;
			LAYER M2 ;
			RECT 17.127 42.680 17.375 42.760 ;
			LAYER M3 ;
			RECT 17.127 42.680 17.375 42.760 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 44.696 17.375 44.776 ;
			LAYER M2 ;
			RECT 17.127 44.696 17.375 44.776 ;
			LAYER M3 ;
			RECT 17.127 44.696 17.375 44.776 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 46.712 17.375 46.792 ;
			LAYER M2 ;
			RECT 17.127 46.712 17.375 46.792 ;
			LAYER M3 ;
			RECT 17.127 46.712 17.375 46.792 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 48.728 17.375 48.808 ;
			LAYER M2 ;
			RECT 17.127 48.728 17.375 48.808 ;
			LAYER M3 ;
			RECT 17.127 48.728 17.375 48.808 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 50.744 17.375 50.824 ;
			LAYER M2 ;
			RECT 17.127 50.744 17.375 50.824 ;
			LAYER M3 ;
			RECT 17.127 50.744 17.375 50.824 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 52.760 17.375 52.840 ;
			LAYER M2 ;
			RECT 17.127 52.760 17.375 52.840 ;
			LAYER M3 ;
			RECT 17.127 52.760 17.375 52.840 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 54.776 17.375 54.856 ;
			LAYER M2 ;
			RECT 17.127 54.776 17.375 54.856 ;
			LAYER M3 ;
			RECT 17.127 54.776 17.375 54.856 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 56.792 17.375 56.872 ;
			LAYER M2 ;
			RECT 17.127 56.792 17.375 56.872 ;
			LAYER M3 ;
			RECT 17.127 56.792 17.375 56.872 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 58.808 17.375 58.888 ;
			LAYER M2 ;
			RECT 17.127 58.808 17.375 58.888 ;
			LAYER M3 ;
			RECT 17.127 58.808 17.375 58.888 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 60.824 17.375 60.904 ;
			LAYER M2 ;
			RECT 17.127 60.824 17.375 60.904 ;
			LAYER M3 ;
			RECT 17.127 60.824 17.375 60.904 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 62.840 17.375 62.920 ;
			LAYER M2 ;
			RECT 17.127 62.840 17.375 62.920 ;
			LAYER M3 ;
			RECT 17.127 62.840 17.375 62.920 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 64.856 17.375 64.936 ;
			LAYER M2 ;
			RECT 17.127 64.856 17.375 64.936 ;
			LAYER M3 ;
			RECT 17.127 64.856 17.375 64.936 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 66.872 17.375 66.952 ;
			LAYER M2 ;
			RECT 17.127 66.872 17.375 66.952 ;
			LAYER M3 ;
			RECT 17.127 66.872 17.375 66.952 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 68.888 17.375 68.968 ;
			LAYER M2 ;
			RECT 17.127 68.888 17.375 68.968 ;
			LAYER M3 ;
			RECT 17.127 68.888 17.375 68.968 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 70.904 17.375 70.984 ;
			LAYER M2 ;
			RECT 17.127 70.904 17.375 70.984 ;
			LAYER M3 ;
			RECT 17.127 70.904 17.375 70.984 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 72.920 17.375 73.000 ;
			LAYER M2 ;
			RECT 17.127 72.920 17.375 73.000 ;
			LAYER M3 ;
			RECT 17.127 72.920 17.375 73.000 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[35]

	PIN D[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 74.936 17.375 75.016 ;
			LAYER M2 ;
			RECT 17.127 74.936 17.375 75.016 ;
			LAYER M3 ;
			RECT 17.127 74.936 17.375 75.016 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[36]

	PIN D[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 76.952 17.375 77.032 ;
			LAYER M2 ;
			RECT 17.127 76.952 17.375 77.032 ;
			LAYER M3 ;
			RECT 17.127 76.952 17.375 77.032 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[37]

	PIN D[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 78.968 17.375 79.048 ;
			LAYER M2 ;
			RECT 17.127 78.968 17.375 79.048 ;
			LAYER M3 ;
			RECT 17.127 78.968 17.375 79.048 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[38]

	PIN D[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 80.984 17.375 81.064 ;
			LAYER M2 ;
			RECT 17.127 80.984 17.375 81.064 ;
			LAYER M3 ;
			RECT 17.127 80.984 17.375 81.064 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[39]

	PIN D[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 83.000 17.375 83.080 ;
			LAYER M2 ;
			RECT 17.127 83.000 17.375 83.080 ;
			LAYER M3 ;
			RECT 17.127 83.000 17.375 83.080 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[40]

	PIN D[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 85.016 17.375 85.096 ;
			LAYER M2 ;
			RECT 17.127 85.016 17.375 85.096 ;
			LAYER M3 ;
			RECT 17.127 85.016 17.375 85.096 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[41]

	PIN D[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 87.032 17.375 87.112 ;
			LAYER M2 ;
			RECT 17.127 87.032 17.375 87.112 ;
			LAYER M3 ;
			RECT 17.127 87.032 17.375 87.112 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[42]

	PIN D[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 89.048 17.375 89.128 ;
			LAYER M2 ;
			RECT 17.127 89.048 17.375 89.128 ;
			LAYER M3 ;
			RECT 17.127 89.048 17.375 89.128 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[43]

	PIN D[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 91.064 17.375 91.144 ;
			LAYER M2 ;
			RECT 17.127 91.064 17.375 91.144 ;
			LAYER M3 ;
			RECT 17.127 91.064 17.375 91.144 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[44]

	PIN D[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 93.080 17.375 93.160 ;
			LAYER M2 ;
			RECT 17.127 93.080 17.375 93.160 ;
			LAYER M3 ;
			RECT 17.127 93.080 17.375 93.160 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[45]

	PIN D[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 95.096 17.375 95.176 ;
			LAYER M2 ;
			RECT 17.127 95.096 17.375 95.176 ;
			LAYER M3 ;
			RECT 17.127 95.096 17.375 95.176 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[46]

	PIN D[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 97.112 17.375 97.192 ;
			LAYER M2 ;
			RECT 17.127 97.112 17.375 97.192 ;
			LAYER M3 ;
			RECT 17.127 97.112 17.375 97.192 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[47]

	PIN D[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 99.128 17.375 99.208 ;
			LAYER M2 ;
			RECT 17.127 99.128 17.375 99.208 ;
			LAYER M3 ;
			RECT 17.127 99.128 17.375 99.208 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[48]

	PIN D[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 101.144 17.375 101.224 ;
			LAYER M2 ;
			RECT 17.127 101.144 17.375 101.224 ;
			LAYER M3 ;
			RECT 17.127 101.144 17.375 101.224 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[49]

	PIN D[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 103.160 17.375 103.240 ;
			LAYER M2 ;
			RECT 17.127 103.160 17.375 103.240 ;
			LAYER M3 ;
			RECT 17.127 103.160 17.375 103.240 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[50]

	PIN D[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 105.176 17.375 105.256 ;
			LAYER M2 ;
			RECT 17.127 105.176 17.375 105.256 ;
			LAYER M3 ;
			RECT 17.127 105.176 17.375 105.256 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[51]

	PIN D[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 107.192 17.375 107.272 ;
			LAYER M2 ;
			RECT 17.127 107.192 17.375 107.272 ;
			LAYER M3 ;
			RECT 17.127 107.192 17.375 107.272 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[52]

	PIN D[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 109.208 17.375 109.288 ;
			LAYER M2 ;
			RECT 17.127 109.208 17.375 109.288 ;
			LAYER M3 ;
			RECT 17.127 109.208 17.375 109.288 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[53]

	PIN D[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 111.224 17.375 111.304 ;
			LAYER M2 ;
			RECT 17.127 111.224 17.375 111.304 ;
			LAYER M3 ;
			RECT 17.127 111.224 17.375 111.304 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[54]

	PIN D[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 113.240 17.375 113.320 ;
			LAYER M2 ;
			RECT 17.127 113.240 17.375 113.320 ;
			LAYER M3 ;
			RECT 17.127 113.240 17.375 113.320 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[55]

	PIN D[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 115.256 17.375 115.336 ;
			LAYER M2 ;
			RECT 17.127 115.256 17.375 115.336 ;
			LAYER M3 ;
			RECT 17.127 115.256 17.375 115.336 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[56]

	PIN D[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 117.272 17.375 117.352 ;
			LAYER M2 ;
			RECT 17.127 117.272 17.375 117.352 ;
			LAYER M3 ;
			RECT 17.127 117.272 17.375 117.352 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[57]

	PIN D[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 119.288 17.375 119.368 ;
			LAYER M2 ;
			RECT 17.127 119.288 17.375 119.368 ;
			LAYER M3 ;
			RECT 17.127 119.288 17.375 119.368 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[58]

	PIN D[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 121.304 17.375 121.384 ;
			LAYER M2 ;
			RECT 17.127 121.304 17.375 121.384 ;
			LAYER M3 ;
			RECT 17.127 121.304 17.375 121.384 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[59]

	PIN D[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 123.320 17.375 123.400 ;
			LAYER M2 ;
			RECT 17.127 123.320 17.375 123.400 ;
			LAYER M3 ;
			RECT 17.127 123.320 17.375 123.400 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[60]

	PIN D[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 125.336 17.375 125.416 ;
			LAYER M2 ;
			RECT 17.127 125.336 17.375 125.416 ;
			LAYER M3 ;
			RECT 17.127 125.336 17.375 125.416 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[61]

	PIN D[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 127.352 17.375 127.432 ;
			LAYER M2 ;
			RECT 17.127 127.352 17.375 127.432 ;
			LAYER M3 ;
			RECT 17.127 127.352 17.375 127.432 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[62]

	PIN D[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 129.368 17.375 129.448 ;
			LAYER M2 ;
			RECT 17.127 129.368 17.375 129.448 ;
			LAYER M3 ;
			RECT 17.127 129.368 17.375 129.448 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[63]

	PIN D[64]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 144.248 17.375 144.328 ;
			LAYER M2 ;
			RECT 17.127 144.248 17.375 144.328 ;
			LAYER M3 ;
			RECT 17.127 144.248 17.375 144.328 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[64]

	PIN D[65]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 146.264 17.375 146.344 ;
			LAYER M2 ;
			RECT 17.127 146.264 17.375 146.344 ;
			LAYER M3 ;
			RECT 17.127 146.264 17.375 146.344 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[65]

	PIN D[66]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 148.280 17.375 148.360 ;
			LAYER M2 ;
			RECT 17.127 148.280 17.375 148.360 ;
			LAYER M3 ;
			RECT 17.127 148.280 17.375 148.360 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[66]

	PIN D[67]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 150.296 17.375 150.376 ;
			LAYER M2 ;
			RECT 17.127 150.296 17.375 150.376 ;
			LAYER M3 ;
			RECT 17.127 150.296 17.375 150.376 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[67]

	PIN D[68]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 152.312 17.375 152.392 ;
			LAYER M2 ;
			RECT 17.127 152.312 17.375 152.392 ;
			LAYER M3 ;
			RECT 17.127 152.312 17.375 152.392 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[68]

	PIN D[69]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 154.328 17.375 154.408 ;
			LAYER M2 ;
			RECT 17.127 154.328 17.375 154.408 ;
			LAYER M3 ;
			RECT 17.127 154.328 17.375 154.408 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[69]

	PIN D[70]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 156.344 17.375 156.424 ;
			LAYER M2 ;
			RECT 17.127 156.344 17.375 156.424 ;
			LAYER M3 ;
			RECT 17.127 156.344 17.375 156.424 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[70]

	PIN D[71]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 158.360 17.375 158.440 ;
			LAYER M2 ;
			RECT 17.127 158.360 17.375 158.440 ;
			LAYER M3 ;
			RECT 17.127 158.360 17.375 158.440 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[71]

	PIN D[72]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 160.376 17.375 160.456 ;
			LAYER M2 ;
			RECT 17.127 160.376 17.375 160.456 ;
			LAYER M3 ;
			RECT 17.127 160.376 17.375 160.456 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[72]

	PIN D[73]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 162.392 17.375 162.472 ;
			LAYER M2 ;
			RECT 17.127 162.392 17.375 162.472 ;
			LAYER M3 ;
			RECT 17.127 162.392 17.375 162.472 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[73]

	PIN D[74]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 164.408 17.375 164.488 ;
			LAYER M2 ;
			RECT 17.127 164.408 17.375 164.488 ;
			LAYER M3 ;
			RECT 17.127 164.408 17.375 164.488 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[74]

	PIN D[75]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 166.424 17.375 166.504 ;
			LAYER M2 ;
			RECT 17.127 166.424 17.375 166.504 ;
			LAYER M3 ;
			RECT 17.127 166.424 17.375 166.504 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[75]

	PIN D[76]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 168.440 17.375 168.520 ;
			LAYER M2 ;
			RECT 17.127 168.440 17.375 168.520 ;
			LAYER M3 ;
			RECT 17.127 168.440 17.375 168.520 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[76]

	PIN D[77]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 170.456 17.375 170.536 ;
			LAYER M2 ;
			RECT 17.127 170.456 17.375 170.536 ;
			LAYER M3 ;
			RECT 17.127 170.456 17.375 170.536 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[77]

	PIN D[78]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 172.472 17.375 172.552 ;
			LAYER M2 ;
			RECT 17.127 172.472 17.375 172.552 ;
			LAYER M3 ;
			RECT 17.127 172.472 17.375 172.552 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[78]

	PIN D[79]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 174.488 17.375 174.568 ;
			LAYER M2 ;
			RECT 17.127 174.488 17.375 174.568 ;
			LAYER M3 ;
			RECT 17.127 174.488 17.375 174.568 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[79]

	PIN D[80]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 176.504 17.375 176.584 ;
			LAYER M2 ;
			RECT 17.127 176.504 17.375 176.584 ;
			LAYER M3 ;
			RECT 17.127 176.504 17.375 176.584 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[80]

	PIN D[81]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 178.520 17.375 178.600 ;
			LAYER M2 ;
			RECT 17.127 178.520 17.375 178.600 ;
			LAYER M3 ;
			RECT 17.127 178.520 17.375 178.600 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[81]

	PIN D[82]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 180.536 17.375 180.616 ;
			LAYER M2 ;
			RECT 17.127 180.536 17.375 180.616 ;
			LAYER M3 ;
			RECT 17.127 180.536 17.375 180.616 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[82]

	PIN D[83]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 182.552 17.375 182.632 ;
			LAYER M2 ;
			RECT 17.127 182.552 17.375 182.632 ;
			LAYER M3 ;
			RECT 17.127 182.552 17.375 182.632 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[83]

	PIN D[84]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 184.568 17.375 184.648 ;
			LAYER M2 ;
			RECT 17.127 184.568 17.375 184.648 ;
			LAYER M3 ;
			RECT 17.127 184.568 17.375 184.648 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[84]

	PIN D[85]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 186.584 17.375 186.664 ;
			LAYER M2 ;
			RECT 17.127 186.584 17.375 186.664 ;
			LAYER M3 ;
			RECT 17.127 186.584 17.375 186.664 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[85]

	PIN D[86]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 188.600 17.375 188.680 ;
			LAYER M2 ;
			RECT 17.127 188.600 17.375 188.680 ;
			LAYER M3 ;
			RECT 17.127 188.600 17.375 188.680 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[86]

	PIN D[87]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 190.616 17.375 190.696 ;
			LAYER M2 ;
			RECT 17.127 190.616 17.375 190.696 ;
			LAYER M3 ;
			RECT 17.127 190.616 17.375 190.696 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[87]

	PIN D[88]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 192.632 17.375 192.712 ;
			LAYER M2 ;
			RECT 17.127 192.632 17.375 192.712 ;
			LAYER M3 ;
			RECT 17.127 192.632 17.375 192.712 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[88]

	PIN D[89]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 194.648 17.375 194.728 ;
			LAYER M2 ;
			RECT 17.127 194.648 17.375 194.728 ;
			LAYER M3 ;
			RECT 17.127 194.648 17.375 194.728 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[89]

	PIN D[90]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 196.664 17.375 196.744 ;
			LAYER M2 ;
			RECT 17.127 196.664 17.375 196.744 ;
			LAYER M3 ;
			RECT 17.127 196.664 17.375 196.744 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[90]

	PIN D[91]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 198.680 17.375 198.760 ;
			LAYER M2 ;
			RECT 17.127 198.680 17.375 198.760 ;
			LAYER M3 ;
			RECT 17.127 198.680 17.375 198.760 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[91]

	PIN D[92]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 200.696 17.375 200.776 ;
			LAYER M2 ;
			RECT 17.127 200.696 17.375 200.776 ;
			LAYER M3 ;
			RECT 17.127 200.696 17.375 200.776 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[92]

	PIN D[93]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 202.712 17.375 202.792 ;
			LAYER M2 ;
			RECT 17.127 202.712 17.375 202.792 ;
			LAYER M3 ;
			RECT 17.127 202.712 17.375 202.792 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[93]

	PIN D[94]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 204.728 17.375 204.808 ;
			LAYER M2 ;
			RECT 17.127 204.728 17.375 204.808 ;
			LAYER M3 ;
			RECT 17.127 204.728 17.375 204.808 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[94]

	PIN D[95]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 206.744 17.375 206.824 ;
			LAYER M2 ;
			RECT 17.127 206.744 17.375 206.824 ;
			LAYER M3 ;
			RECT 17.127 206.744 17.375 206.824 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[95]

	PIN D[96]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 208.760 17.375 208.840 ;
			LAYER M2 ;
			RECT 17.127 208.760 17.375 208.840 ;
			LAYER M3 ;
			RECT 17.127 208.760 17.375 208.840 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[96]

	PIN D[97]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 210.776 17.375 210.856 ;
			LAYER M2 ;
			RECT 17.127 210.776 17.375 210.856 ;
			LAYER M3 ;
			RECT 17.127 210.776 17.375 210.856 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[97]

	PIN D[98]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 212.792 17.375 212.872 ;
			LAYER M2 ;
			RECT 17.127 212.792 17.375 212.872 ;
			LAYER M3 ;
			RECT 17.127 212.792 17.375 212.872 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[98]

	PIN D[99]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 214.808 17.375 214.888 ;
			LAYER M2 ;
			RECT 17.127 214.808 17.375 214.888 ;
			LAYER M3 ;
			RECT 17.127 214.808 17.375 214.888 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[99]

	PIN D[100]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 216.824 17.375 216.904 ;
			LAYER M2 ;
			RECT 17.127 216.824 17.375 216.904 ;
			LAYER M3 ;
			RECT 17.127 216.824 17.375 216.904 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[100]

	PIN D[101]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 218.840 17.375 218.920 ;
			LAYER M2 ;
			RECT 17.127 218.840 17.375 218.920 ;
			LAYER M3 ;
			RECT 17.127 218.840 17.375 218.920 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[101]

	PIN D[102]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 220.856 17.375 220.936 ;
			LAYER M2 ;
			RECT 17.127 220.856 17.375 220.936 ;
			LAYER M3 ;
			RECT 17.127 220.856 17.375 220.936 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[102]

	PIN D[103]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 222.872 17.375 222.952 ;
			LAYER M2 ;
			RECT 17.127 222.872 17.375 222.952 ;
			LAYER M3 ;
			RECT 17.127 222.872 17.375 222.952 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[103]

	PIN D[104]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 224.888 17.375 224.968 ;
			LAYER M2 ;
			RECT 17.127 224.888 17.375 224.968 ;
			LAYER M3 ;
			RECT 17.127 224.888 17.375 224.968 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[104]

	PIN D[105]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 226.904 17.375 226.984 ;
			LAYER M2 ;
			RECT 17.127 226.904 17.375 226.984 ;
			LAYER M3 ;
			RECT 17.127 226.904 17.375 226.984 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[105]

	PIN D[106]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 228.920 17.375 229.000 ;
			LAYER M2 ;
			RECT 17.127 228.920 17.375 229.000 ;
			LAYER M3 ;
			RECT 17.127 228.920 17.375 229.000 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[106]

	PIN D[107]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 230.936 17.375 231.016 ;
			LAYER M2 ;
			RECT 17.127 230.936 17.375 231.016 ;
			LAYER M3 ;
			RECT 17.127 230.936 17.375 231.016 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[107]

	PIN D[108]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 232.952 17.375 233.032 ;
			LAYER M2 ;
			RECT 17.127 232.952 17.375 233.032 ;
			LAYER M3 ;
			RECT 17.127 232.952 17.375 233.032 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[108]

	PIN D[109]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 234.968 17.375 235.048 ;
			LAYER M2 ;
			RECT 17.127 234.968 17.375 235.048 ;
			LAYER M3 ;
			RECT 17.127 234.968 17.375 235.048 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[109]

	PIN D[110]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 236.984 17.375 237.064 ;
			LAYER M2 ;
			RECT 17.127 236.984 17.375 237.064 ;
			LAYER M3 ;
			RECT 17.127 236.984 17.375 237.064 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[110]

	PIN D[111]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 239.000 17.375 239.080 ;
			LAYER M2 ;
			RECT 17.127 239.000 17.375 239.080 ;
			LAYER M3 ;
			RECT 17.127 239.000 17.375 239.080 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[111]

	PIN D[112]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 241.016 17.375 241.096 ;
			LAYER M2 ;
			RECT 17.127 241.016 17.375 241.096 ;
			LAYER M3 ;
			RECT 17.127 241.016 17.375 241.096 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[112]

	PIN D[113]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 243.032 17.375 243.112 ;
			LAYER M2 ;
			RECT 17.127 243.032 17.375 243.112 ;
			LAYER M3 ;
			RECT 17.127 243.032 17.375 243.112 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[113]

	PIN D[114]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 245.048 17.375 245.128 ;
			LAYER M2 ;
			RECT 17.127 245.048 17.375 245.128 ;
			LAYER M3 ;
			RECT 17.127 245.048 17.375 245.128 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[114]

	PIN D[115]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 247.064 17.375 247.144 ;
			LAYER M2 ;
			RECT 17.127 247.064 17.375 247.144 ;
			LAYER M3 ;
			RECT 17.127 247.064 17.375 247.144 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[115]

	PIN D[116]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 249.080 17.375 249.160 ;
			LAYER M2 ;
			RECT 17.127 249.080 17.375 249.160 ;
			LAYER M3 ;
			RECT 17.127 249.080 17.375 249.160 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[116]

	PIN D[117]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 251.096 17.375 251.176 ;
			LAYER M2 ;
			RECT 17.127 251.096 17.375 251.176 ;
			LAYER M3 ;
			RECT 17.127 251.096 17.375 251.176 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[117]

	PIN D[118]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 253.112 17.375 253.192 ;
			LAYER M2 ;
			RECT 17.127 253.112 17.375 253.192 ;
			LAYER M3 ;
			RECT 17.127 253.112 17.375 253.192 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[118]

	PIN D[119]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 255.128 17.375 255.208 ;
			LAYER M2 ;
			RECT 17.127 255.128 17.375 255.208 ;
			LAYER M3 ;
			RECT 17.127 255.128 17.375 255.208 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[119]

	PIN D[120]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 257.144 17.375 257.224 ;
			LAYER M2 ;
			RECT 17.127 257.144 17.375 257.224 ;
			LAYER M3 ;
			RECT 17.127 257.144 17.375 257.224 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[120]

	PIN D[121]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 259.160 17.375 259.240 ;
			LAYER M2 ;
			RECT 17.127 259.160 17.375 259.240 ;
			LAYER M3 ;
			RECT 17.127 259.160 17.375 259.240 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[121]

	PIN D[122]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 261.176 17.375 261.256 ;
			LAYER M2 ;
			RECT 17.127 261.176 17.375 261.256 ;
			LAYER M3 ;
			RECT 17.127 261.176 17.375 261.256 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[122]

	PIN D[123]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 263.192 17.375 263.272 ;
			LAYER M2 ;
			RECT 17.127 263.192 17.375 263.272 ;
			LAYER M3 ;
			RECT 17.127 263.192 17.375 263.272 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[123]

	PIN D[124]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 265.208 17.375 265.288 ;
			LAYER M2 ;
			RECT 17.127 265.208 17.375 265.288 ;
			LAYER M3 ;
			RECT 17.127 265.208 17.375 265.288 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[124]

	PIN D[125]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 267.224 17.375 267.304 ;
			LAYER M2 ;
			RECT 17.127 267.224 17.375 267.304 ;
			LAYER M3 ;
			RECT 17.127 267.224 17.375 267.304 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[125]

	PIN D[126]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 269.240 17.375 269.320 ;
			LAYER M2 ;
			RECT 17.127 269.240 17.375 269.320 ;
			LAYER M3 ;
			RECT 17.127 269.240 17.375 269.320 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[126]

	PIN D[127]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 271.256 17.375 271.336 ;
			LAYER M2 ;
			RECT 17.127 271.256 17.375 271.336 ;
			LAYER M3 ;
			RECT 17.127 271.256 17.375 271.336 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[127]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 1.208 17.375 1.288 ;
			LAYER M2 ;
			RECT 17.127 1.208 17.375 1.288 ;
			LAYER M3 ;
			RECT 17.127 1.208 17.375 1.288 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 3.224 17.375 3.304 ;
			LAYER M2 ;
			RECT 17.127 3.224 17.375 3.304 ;
			LAYER M3 ;
			RECT 17.127 3.224 17.375 3.304 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 5.240 17.375 5.320 ;
			LAYER M2 ;
			RECT 17.127 5.240 17.375 5.320 ;
			LAYER M3 ;
			RECT 17.127 5.240 17.375 5.320 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 7.256 17.375 7.336 ;
			LAYER M2 ;
			RECT 17.127 7.256 17.375 7.336 ;
			LAYER M3 ;
			RECT 17.127 7.256 17.375 7.336 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 9.272 17.375 9.352 ;
			LAYER M2 ;
			RECT 17.127 9.272 17.375 9.352 ;
			LAYER M3 ;
			RECT 17.127 9.272 17.375 9.352 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 11.288 17.375 11.368 ;
			LAYER M2 ;
			RECT 17.127 11.288 17.375 11.368 ;
			LAYER M3 ;
			RECT 17.127 11.288 17.375 11.368 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 13.304 17.375 13.384 ;
			LAYER M2 ;
			RECT 17.127 13.304 17.375 13.384 ;
			LAYER M3 ;
			RECT 17.127 13.304 17.375 13.384 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 15.320 17.375 15.400 ;
			LAYER M2 ;
			RECT 17.127 15.320 17.375 15.400 ;
			LAYER M3 ;
			RECT 17.127 15.320 17.375 15.400 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 17.336 17.375 17.416 ;
			LAYER M2 ;
			RECT 17.127 17.336 17.375 17.416 ;
			LAYER M3 ;
			RECT 17.127 17.336 17.375 17.416 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 19.352 17.375 19.432 ;
			LAYER M2 ;
			RECT 17.127 19.352 17.375 19.432 ;
			LAYER M3 ;
			RECT 17.127 19.352 17.375 19.432 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 21.368 17.375 21.448 ;
			LAYER M2 ;
			RECT 17.127 21.368 17.375 21.448 ;
			LAYER M3 ;
			RECT 17.127 21.368 17.375 21.448 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 23.384 17.375 23.464 ;
			LAYER M2 ;
			RECT 17.127 23.384 17.375 23.464 ;
			LAYER M3 ;
			RECT 17.127 23.384 17.375 23.464 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 25.400 17.375 25.480 ;
			LAYER M2 ;
			RECT 17.127 25.400 17.375 25.480 ;
			LAYER M3 ;
			RECT 17.127 25.400 17.375 25.480 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 27.416 17.375 27.496 ;
			LAYER M2 ;
			RECT 17.127 27.416 17.375 27.496 ;
			LAYER M3 ;
			RECT 17.127 27.416 17.375 27.496 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 29.432 17.375 29.512 ;
			LAYER M2 ;
			RECT 17.127 29.432 17.375 29.512 ;
			LAYER M3 ;
			RECT 17.127 29.432 17.375 29.512 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 31.448 17.375 31.528 ;
			LAYER M2 ;
			RECT 17.127 31.448 17.375 31.528 ;
			LAYER M3 ;
			RECT 17.127 31.448 17.375 31.528 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 33.464 17.375 33.544 ;
			LAYER M2 ;
			RECT 17.127 33.464 17.375 33.544 ;
			LAYER M3 ;
			RECT 17.127 33.464 17.375 33.544 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 35.480 17.375 35.560 ;
			LAYER M2 ;
			RECT 17.127 35.480 17.375 35.560 ;
			LAYER M3 ;
			RECT 17.127 35.480 17.375 35.560 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 37.496 17.375 37.576 ;
			LAYER M2 ;
			RECT 17.127 37.496 17.375 37.576 ;
			LAYER M3 ;
			RECT 17.127 37.496 17.375 37.576 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 39.512 17.375 39.592 ;
			LAYER M2 ;
			RECT 17.127 39.512 17.375 39.592 ;
			LAYER M3 ;
			RECT 17.127 39.512 17.375 39.592 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 41.528 17.375 41.608 ;
			LAYER M2 ;
			RECT 17.127 41.528 17.375 41.608 ;
			LAYER M3 ;
			RECT 17.127 41.528 17.375 41.608 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 43.544 17.375 43.624 ;
			LAYER M2 ;
			RECT 17.127 43.544 17.375 43.624 ;
			LAYER M3 ;
			RECT 17.127 43.544 17.375 43.624 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 45.560 17.375 45.640 ;
			LAYER M2 ;
			RECT 17.127 45.560 17.375 45.640 ;
			LAYER M3 ;
			RECT 17.127 45.560 17.375 45.640 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 47.576 17.375 47.656 ;
			LAYER M2 ;
			RECT 17.127 47.576 17.375 47.656 ;
			LAYER M3 ;
			RECT 17.127 47.576 17.375 47.656 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 49.592 17.375 49.672 ;
			LAYER M2 ;
			RECT 17.127 49.592 17.375 49.672 ;
			LAYER M3 ;
			RECT 17.127 49.592 17.375 49.672 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 51.608 17.375 51.688 ;
			LAYER M2 ;
			RECT 17.127 51.608 17.375 51.688 ;
			LAYER M3 ;
			RECT 17.127 51.608 17.375 51.688 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 53.624 17.375 53.704 ;
			LAYER M2 ;
			RECT 17.127 53.624 17.375 53.704 ;
			LAYER M3 ;
			RECT 17.127 53.624 17.375 53.704 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 55.640 17.375 55.720 ;
			LAYER M2 ;
			RECT 17.127 55.640 17.375 55.720 ;
			LAYER M3 ;
			RECT 17.127 55.640 17.375 55.720 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 57.656 17.375 57.736 ;
			LAYER M2 ;
			RECT 17.127 57.656 17.375 57.736 ;
			LAYER M3 ;
			RECT 17.127 57.656 17.375 57.736 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 59.672 17.375 59.752 ;
			LAYER M2 ;
			RECT 17.127 59.672 17.375 59.752 ;
			LAYER M3 ;
			RECT 17.127 59.672 17.375 59.752 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 61.688 17.375 61.768 ;
			LAYER M2 ;
			RECT 17.127 61.688 17.375 61.768 ;
			LAYER M3 ;
			RECT 17.127 61.688 17.375 61.768 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 63.704 17.375 63.784 ;
			LAYER M2 ;
			RECT 17.127 63.704 17.375 63.784 ;
			LAYER M3 ;
			RECT 17.127 63.704 17.375 63.784 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 65.720 17.375 65.800 ;
			LAYER M2 ;
			RECT 17.127 65.720 17.375 65.800 ;
			LAYER M3 ;
			RECT 17.127 65.720 17.375 65.800 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 67.736 17.375 67.816 ;
			LAYER M2 ;
			RECT 17.127 67.736 17.375 67.816 ;
			LAYER M3 ;
			RECT 17.127 67.736 17.375 67.816 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 69.752 17.375 69.832 ;
			LAYER M2 ;
			RECT 17.127 69.752 17.375 69.832 ;
			LAYER M3 ;
			RECT 17.127 69.752 17.375 69.832 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 71.768 17.375 71.848 ;
			LAYER M2 ;
			RECT 17.127 71.768 17.375 71.848 ;
			LAYER M3 ;
			RECT 17.127 71.768 17.375 71.848 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[35]

	PIN Q[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 73.784 17.375 73.864 ;
			LAYER M2 ;
			RECT 17.127 73.784 17.375 73.864 ;
			LAYER M3 ;
			RECT 17.127 73.784 17.375 73.864 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[36]

	PIN Q[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 75.800 17.375 75.880 ;
			LAYER M2 ;
			RECT 17.127 75.800 17.375 75.880 ;
			LAYER M3 ;
			RECT 17.127 75.800 17.375 75.880 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[37]

	PIN Q[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 77.816 17.375 77.896 ;
			LAYER M2 ;
			RECT 17.127 77.816 17.375 77.896 ;
			LAYER M3 ;
			RECT 17.127 77.816 17.375 77.896 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[38]

	PIN Q[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 79.832 17.375 79.912 ;
			LAYER M2 ;
			RECT 17.127 79.832 17.375 79.912 ;
			LAYER M3 ;
			RECT 17.127 79.832 17.375 79.912 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[39]

	PIN Q[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 81.848 17.375 81.928 ;
			LAYER M2 ;
			RECT 17.127 81.848 17.375 81.928 ;
			LAYER M3 ;
			RECT 17.127 81.848 17.375 81.928 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[40]

	PIN Q[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 83.864 17.375 83.944 ;
			LAYER M2 ;
			RECT 17.127 83.864 17.375 83.944 ;
			LAYER M3 ;
			RECT 17.127 83.864 17.375 83.944 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[41]

	PIN Q[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 85.880 17.375 85.960 ;
			LAYER M2 ;
			RECT 17.127 85.880 17.375 85.960 ;
			LAYER M3 ;
			RECT 17.127 85.880 17.375 85.960 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[42]

	PIN Q[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 87.896 17.375 87.976 ;
			LAYER M2 ;
			RECT 17.127 87.896 17.375 87.976 ;
			LAYER M3 ;
			RECT 17.127 87.896 17.375 87.976 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[43]

	PIN Q[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 89.912 17.375 89.992 ;
			LAYER M2 ;
			RECT 17.127 89.912 17.375 89.992 ;
			LAYER M3 ;
			RECT 17.127 89.912 17.375 89.992 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[44]

	PIN Q[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 91.928 17.375 92.008 ;
			LAYER M2 ;
			RECT 17.127 91.928 17.375 92.008 ;
			LAYER M3 ;
			RECT 17.127 91.928 17.375 92.008 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[45]

	PIN Q[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 93.944 17.375 94.024 ;
			LAYER M2 ;
			RECT 17.127 93.944 17.375 94.024 ;
			LAYER M3 ;
			RECT 17.127 93.944 17.375 94.024 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[46]

	PIN Q[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 95.960 17.375 96.040 ;
			LAYER M2 ;
			RECT 17.127 95.960 17.375 96.040 ;
			LAYER M3 ;
			RECT 17.127 95.960 17.375 96.040 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[47]

	PIN Q[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 97.976 17.375 98.056 ;
			LAYER M2 ;
			RECT 17.127 97.976 17.375 98.056 ;
			LAYER M3 ;
			RECT 17.127 97.976 17.375 98.056 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[48]

	PIN Q[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 99.992 17.375 100.072 ;
			LAYER M2 ;
			RECT 17.127 99.992 17.375 100.072 ;
			LAYER M3 ;
			RECT 17.127 99.992 17.375 100.072 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[49]

	PIN Q[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 102.008 17.375 102.088 ;
			LAYER M2 ;
			RECT 17.127 102.008 17.375 102.088 ;
			LAYER M3 ;
			RECT 17.127 102.008 17.375 102.088 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[50]

	PIN Q[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 104.024 17.375 104.104 ;
			LAYER M2 ;
			RECT 17.127 104.024 17.375 104.104 ;
			LAYER M3 ;
			RECT 17.127 104.024 17.375 104.104 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[51]

	PIN Q[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 106.040 17.375 106.120 ;
			LAYER M2 ;
			RECT 17.127 106.040 17.375 106.120 ;
			LAYER M3 ;
			RECT 17.127 106.040 17.375 106.120 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[52]

	PIN Q[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 108.056 17.375 108.136 ;
			LAYER M2 ;
			RECT 17.127 108.056 17.375 108.136 ;
			LAYER M3 ;
			RECT 17.127 108.056 17.375 108.136 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[53]

	PIN Q[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 110.072 17.375 110.152 ;
			LAYER M2 ;
			RECT 17.127 110.072 17.375 110.152 ;
			LAYER M3 ;
			RECT 17.127 110.072 17.375 110.152 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[54]

	PIN Q[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 112.088 17.375 112.168 ;
			LAYER M2 ;
			RECT 17.127 112.088 17.375 112.168 ;
			LAYER M3 ;
			RECT 17.127 112.088 17.375 112.168 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[55]

	PIN Q[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 114.104 17.375 114.184 ;
			LAYER M2 ;
			RECT 17.127 114.104 17.375 114.184 ;
			LAYER M3 ;
			RECT 17.127 114.104 17.375 114.184 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[56]

	PIN Q[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 116.120 17.375 116.200 ;
			LAYER M2 ;
			RECT 17.127 116.120 17.375 116.200 ;
			LAYER M3 ;
			RECT 17.127 116.120 17.375 116.200 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[57]

	PIN Q[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 118.136 17.375 118.216 ;
			LAYER M2 ;
			RECT 17.127 118.136 17.375 118.216 ;
			LAYER M3 ;
			RECT 17.127 118.136 17.375 118.216 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[58]

	PIN Q[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 120.152 17.375 120.232 ;
			LAYER M2 ;
			RECT 17.127 120.152 17.375 120.232 ;
			LAYER M3 ;
			RECT 17.127 120.152 17.375 120.232 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[59]

	PIN Q[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 122.168 17.375 122.248 ;
			LAYER M2 ;
			RECT 17.127 122.168 17.375 122.248 ;
			LAYER M3 ;
			RECT 17.127 122.168 17.375 122.248 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[60]

	PIN Q[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 124.184 17.375 124.264 ;
			LAYER M2 ;
			RECT 17.127 124.184 17.375 124.264 ;
			LAYER M3 ;
			RECT 17.127 124.184 17.375 124.264 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[61]

	PIN Q[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 126.200 17.375 126.280 ;
			LAYER M2 ;
			RECT 17.127 126.200 17.375 126.280 ;
			LAYER M3 ;
			RECT 17.127 126.200 17.375 126.280 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[62]

	PIN Q[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 128.216 17.375 128.296 ;
			LAYER M2 ;
			RECT 17.127 128.216 17.375 128.296 ;
			LAYER M3 ;
			RECT 17.127 128.216 17.375 128.296 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[63]

	PIN Q[64]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 143.096 17.375 143.176 ;
			LAYER M2 ;
			RECT 17.127 143.096 17.375 143.176 ;
			LAYER M3 ;
			RECT 17.127 143.096 17.375 143.176 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[64]

	PIN Q[65]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 145.112 17.375 145.192 ;
			LAYER M2 ;
			RECT 17.127 145.112 17.375 145.192 ;
			LAYER M3 ;
			RECT 17.127 145.112 17.375 145.192 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[65]

	PIN Q[66]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 147.128 17.375 147.208 ;
			LAYER M2 ;
			RECT 17.127 147.128 17.375 147.208 ;
			LAYER M3 ;
			RECT 17.127 147.128 17.375 147.208 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[66]

	PIN Q[67]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 149.144 17.375 149.224 ;
			LAYER M2 ;
			RECT 17.127 149.144 17.375 149.224 ;
			LAYER M3 ;
			RECT 17.127 149.144 17.375 149.224 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[67]

	PIN Q[68]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 151.160 17.375 151.240 ;
			LAYER M2 ;
			RECT 17.127 151.160 17.375 151.240 ;
			LAYER M3 ;
			RECT 17.127 151.160 17.375 151.240 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[68]

	PIN Q[69]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 153.176 17.375 153.256 ;
			LAYER M2 ;
			RECT 17.127 153.176 17.375 153.256 ;
			LAYER M3 ;
			RECT 17.127 153.176 17.375 153.256 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[69]

	PIN Q[70]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 155.192 17.375 155.272 ;
			LAYER M2 ;
			RECT 17.127 155.192 17.375 155.272 ;
			LAYER M3 ;
			RECT 17.127 155.192 17.375 155.272 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[70]

	PIN Q[71]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 157.208 17.375 157.288 ;
			LAYER M2 ;
			RECT 17.127 157.208 17.375 157.288 ;
			LAYER M3 ;
			RECT 17.127 157.208 17.375 157.288 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[71]

	PIN Q[72]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 159.224 17.375 159.304 ;
			LAYER M2 ;
			RECT 17.127 159.224 17.375 159.304 ;
			LAYER M3 ;
			RECT 17.127 159.224 17.375 159.304 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[72]

	PIN Q[73]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 161.240 17.375 161.320 ;
			LAYER M2 ;
			RECT 17.127 161.240 17.375 161.320 ;
			LAYER M3 ;
			RECT 17.127 161.240 17.375 161.320 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[73]

	PIN Q[74]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 163.256 17.375 163.336 ;
			LAYER M2 ;
			RECT 17.127 163.256 17.375 163.336 ;
			LAYER M3 ;
			RECT 17.127 163.256 17.375 163.336 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[74]

	PIN Q[75]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 165.272 17.375 165.352 ;
			LAYER M2 ;
			RECT 17.127 165.272 17.375 165.352 ;
			LAYER M3 ;
			RECT 17.127 165.272 17.375 165.352 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[75]

	PIN Q[76]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 167.288 17.375 167.368 ;
			LAYER M2 ;
			RECT 17.127 167.288 17.375 167.368 ;
			LAYER M3 ;
			RECT 17.127 167.288 17.375 167.368 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[76]

	PIN Q[77]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 169.304 17.375 169.384 ;
			LAYER M2 ;
			RECT 17.127 169.304 17.375 169.384 ;
			LAYER M3 ;
			RECT 17.127 169.304 17.375 169.384 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[77]

	PIN Q[78]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 171.320 17.375 171.400 ;
			LAYER M2 ;
			RECT 17.127 171.320 17.375 171.400 ;
			LAYER M3 ;
			RECT 17.127 171.320 17.375 171.400 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[78]

	PIN Q[79]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 173.336 17.375 173.416 ;
			LAYER M2 ;
			RECT 17.127 173.336 17.375 173.416 ;
			LAYER M3 ;
			RECT 17.127 173.336 17.375 173.416 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[79]

	PIN Q[80]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 175.352 17.375 175.432 ;
			LAYER M2 ;
			RECT 17.127 175.352 17.375 175.432 ;
			LAYER M3 ;
			RECT 17.127 175.352 17.375 175.432 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[80]

	PIN Q[81]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 177.368 17.375 177.448 ;
			LAYER M2 ;
			RECT 17.127 177.368 17.375 177.448 ;
			LAYER M3 ;
			RECT 17.127 177.368 17.375 177.448 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[81]

	PIN Q[82]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 179.384 17.375 179.464 ;
			LAYER M2 ;
			RECT 17.127 179.384 17.375 179.464 ;
			LAYER M3 ;
			RECT 17.127 179.384 17.375 179.464 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[82]

	PIN Q[83]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 181.400 17.375 181.480 ;
			LAYER M2 ;
			RECT 17.127 181.400 17.375 181.480 ;
			LAYER M3 ;
			RECT 17.127 181.400 17.375 181.480 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[83]

	PIN Q[84]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 183.416 17.375 183.496 ;
			LAYER M2 ;
			RECT 17.127 183.416 17.375 183.496 ;
			LAYER M3 ;
			RECT 17.127 183.416 17.375 183.496 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[84]

	PIN Q[85]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 185.432 17.375 185.512 ;
			LAYER M2 ;
			RECT 17.127 185.432 17.375 185.512 ;
			LAYER M3 ;
			RECT 17.127 185.432 17.375 185.512 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[85]

	PIN Q[86]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 187.448 17.375 187.528 ;
			LAYER M2 ;
			RECT 17.127 187.448 17.375 187.528 ;
			LAYER M3 ;
			RECT 17.127 187.448 17.375 187.528 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[86]

	PIN Q[87]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 189.464 17.375 189.544 ;
			LAYER M2 ;
			RECT 17.127 189.464 17.375 189.544 ;
			LAYER M3 ;
			RECT 17.127 189.464 17.375 189.544 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[87]

	PIN Q[88]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 191.480 17.375 191.560 ;
			LAYER M2 ;
			RECT 17.127 191.480 17.375 191.560 ;
			LAYER M3 ;
			RECT 17.127 191.480 17.375 191.560 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[88]

	PIN Q[89]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 193.496 17.375 193.576 ;
			LAYER M2 ;
			RECT 17.127 193.496 17.375 193.576 ;
			LAYER M3 ;
			RECT 17.127 193.496 17.375 193.576 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[89]

	PIN Q[90]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 195.512 17.375 195.592 ;
			LAYER M2 ;
			RECT 17.127 195.512 17.375 195.592 ;
			LAYER M3 ;
			RECT 17.127 195.512 17.375 195.592 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[90]

	PIN Q[91]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 197.528 17.375 197.608 ;
			LAYER M2 ;
			RECT 17.127 197.528 17.375 197.608 ;
			LAYER M3 ;
			RECT 17.127 197.528 17.375 197.608 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[91]

	PIN Q[92]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 199.544 17.375 199.624 ;
			LAYER M2 ;
			RECT 17.127 199.544 17.375 199.624 ;
			LAYER M3 ;
			RECT 17.127 199.544 17.375 199.624 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[92]

	PIN Q[93]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 201.560 17.375 201.640 ;
			LAYER M2 ;
			RECT 17.127 201.560 17.375 201.640 ;
			LAYER M3 ;
			RECT 17.127 201.560 17.375 201.640 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[93]

	PIN Q[94]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 203.576 17.375 203.656 ;
			LAYER M2 ;
			RECT 17.127 203.576 17.375 203.656 ;
			LAYER M3 ;
			RECT 17.127 203.576 17.375 203.656 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[94]

	PIN Q[95]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 205.592 17.375 205.672 ;
			LAYER M2 ;
			RECT 17.127 205.592 17.375 205.672 ;
			LAYER M3 ;
			RECT 17.127 205.592 17.375 205.672 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[95]

	PIN Q[96]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 207.608 17.375 207.688 ;
			LAYER M2 ;
			RECT 17.127 207.608 17.375 207.688 ;
			LAYER M3 ;
			RECT 17.127 207.608 17.375 207.688 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[96]

	PIN Q[97]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 209.624 17.375 209.704 ;
			LAYER M2 ;
			RECT 17.127 209.624 17.375 209.704 ;
			LAYER M3 ;
			RECT 17.127 209.624 17.375 209.704 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[97]

	PIN Q[98]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 211.640 17.375 211.720 ;
			LAYER M2 ;
			RECT 17.127 211.640 17.375 211.720 ;
			LAYER M3 ;
			RECT 17.127 211.640 17.375 211.720 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[98]

	PIN Q[99]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 213.656 17.375 213.736 ;
			LAYER M2 ;
			RECT 17.127 213.656 17.375 213.736 ;
			LAYER M3 ;
			RECT 17.127 213.656 17.375 213.736 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[99]

	PIN Q[100]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 215.672 17.375 215.752 ;
			LAYER M2 ;
			RECT 17.127 215.672 17.375 215.752 ;
			LAYER M3 ;
			RECT 17.127 215.672 17.375 215.752 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[100]

	PIN Q[101]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 217.688 17.375 217.768 ;
			LAYER M2 ;
			RECT 17.127 217.688 17.375 217.768 ;
			LAYER M3 ;
			RECT 17.127 217.688 17.375 217.768 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[101]

	PIN Q[102]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 219.704 17.375 219.784 ;
			LAYER M2 ;
			RECT 17.127 219.704 17.375 219.784 ;
			LAYER M3 ;
			RECT 17.127 219.704 17.375 219.784 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[102]

	PIN Q[103]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 221.720 17.375 221.800 ;
			LAYER M2 ;
			RECT 17.127 221.720 17.375 221.800 ;
			LAYER M3 ;
			RECT 17.127 221.720 17.375 221.800 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[103]

	PIN Q[104]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 223.736 17.375 223.816 ;
			LAYER M2 ;
			RECT 17.127 223.736 17.375 223.816 ;
			LAYER M3 ;
			RECT 17.127 223.736 17.375 223.816 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[104]

	PIN Q[105]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 225.752 17.375 225.832 ;
			LAYER M2 ;
			RECT 17.127 225.752 17.375 225.832 ;
			LAYER M3 ;
			RECT 17.127 225.752 17.375 225.832 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[105]

	PIN Q[106]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 227.768 17.375 227.848 ;
			LAYER M2 ;
			RECT 17.127 227.768 17.375 227.848 ;
			LAYER M3 ;
			RECT 17.127 227.768 17.375 227.848 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[106]

	PIN Q[107]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 229.784 17.375 229.864 ;
			LAYER M2 ;
			RECT 17.127 229.784 17.375 229.864 ;
			LAYER M3 ;
			RECT 17.127 229.784 17.375 229.864 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[107]

	PIN Q[108]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 231.800 17.375 231.880 ;
			LAYER M2 ;
			RECT 17.127 231.800 17.375 231.880 ;
			LAYER M3 ;
			RECT 17.127 231.800 17.375 231.880 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[108]

	PIN Q[109]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 233.816 17.375 233.896 ;
			LAYER M2 ;
			RECT 17.127 233.816 17.375 233.896 ;
			LAYER M3 ;
			RECT 17.127 233.816 17.375 233.896 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[109]

	PIN Q[110]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 235.832 17.375 235.912 ;
			LAYER M2 ;
			RECT 17.127 235.832 17.375 235.912 ;
			LAYER M3 ;
			RECT 17.127 235.832 17.375 235.912 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[110]

	PIN Q[111]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 237.848 17.375 237.928 ;
			LAYER M2 ;
			RECT 17.127 237.848 17.375 237.928 ;
			LAYER M3 ;
			RECT 17.127 237.848 17.375 237.928 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[111]

	PIN Q[112]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 239.864 17.375 239.944 ;
			LAYER M2 ;
			RECT 17.127 239.864 17.375 239.944 ;
			LAYER M3 ;
			RECT 17.127 239.864 17.375 239.944 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[112]

	PIN Q[113]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 241.880 17.375 241.960 ;
			LAYER M2 ;
			RECT 17.127 241.880 17.375 241.960 ;
			LAYER M3 ;
			RECT 17.127 241.880 17.375 241.960 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[113]

	PIN Q[114]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 243.896 17.375 243.976 ;
			LAYER M2 ;
			RECT 17.127 243.896 17.375 243.976 ;
			LAYER M3 ;
			RECT 17.127 243.896 17.375 243.976 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[114]

	PIN Q[115]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 245.912 17.375 245.992 ;
			LAYER M2 ;
			RECT 17.127 245.912 17.375 245.992 ;
			LAYER M3 ;
			RECT 17.127 245.912 17.375 245.992 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[115]

	PIN Q[116]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 247.928 17.375 248.008 ;
			LAYER M2 ;
			RECT 17.127 247.928 17.375 248.008 ;
			LAYER M3 ;
			RECT 17.127 247.928 17.375 248.008 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[116]

	PIN Q[117]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 249.944 17.375 250.024 ;
			LAYER M2 ;
			RECT 17.127 249.944 17.375 250.024 ;
			LAYER M3 ;
			RECT 17.127 249.944 17.375 250.024 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[117]

	PIN Q[118]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 251.960 17.375 252.040 ;
			LAYER M2 ;
			RECT 17.127 251.960 17.375 252.040 ;
			LAYER M3 ;
			RECT 17.127 251.960 17.375 252.040 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[118]

	PIN Q[119]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 253.976 17.375 254.056 ;
			LAYER M2 ;
			RECT 17.127 253.976 17.375 254.056 ;
			LAYER M3 ;
			RECT 17.127 253.976 17.375 254.056 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[119]

	PIN Q[120]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 255.992 17.375 256.072 ;
			LAYER M2 ;
			RECT 17.127 255.992 17.375 256.072 ;
			LAYER M3 ;
			RECT 17.127 255.992 17.375 256.072 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[120]

	PIN Q[121]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 258.008 17.375 258.088 ;
			LAYER M2 ;
			RECT 17.127 258.008 17.375 258.088 ;
			LAYER M3 ;
			RECT 17.127 258.008 17.375 258.088 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[121]

	PIN Q[122]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 260.024 17.375 260.104 ;
			LAYER M2 ;
			RECT 17.127 260.024 17.375 260.104 ;
			LAYER M3 ;
			RECT 17.127 260.024 17.375 260.104 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[122]

	PIN Q[123]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 262.040 17.375 262.120 ;
			LAYER M2 ;
			RECT 17.127 262.040 17.375 262.120 ;
			LAYER M3 ;
			RECT 17.127 262.040 17.375 262.120 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[123]

	PIN Q[124]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 264.056 17.375 264.136 ;
			LAYER M2 ;
			RECT 17.127 264.056 17.375 264.136 ;
			LAYER M3 ;
			RECT 17.127 264.056 17.375 264.136 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[124]

	PIN Q[125]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 266.072 17.375 266.152 ;
			LAYER M2 ;
			RECT 17.127 266.072 17.375 266.152 ;
			LAYER M3 ;
			RECT 17.127 266.072 17.375 266.152 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[125]

	PIN Q[126]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 268.088 17.375 268.168 ;
			LAYER M2 ;
			RECT 17.127 268.088 17.375 268.168 ;
			LAYER M3 ;
			RECT 17.127 268.088 17.375 268.168 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[126]

	PIN Q[127]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 270.104 17.375 270.184 ;
			LAYER M2 ;
			RECT 17.127 270.104 17.375 270.184 ;
			LAYER M3 ;
			RECT 17.127 270.104 17.375 270.184 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[127]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 141.704 17.375 141.784 ;
			LAYER M2 ;
			RECT 17.127 141.704 17.375 141.784 ;
			LAYER M3 ;
			RECT 17.127 141.704 17.375 141.784 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128800 LAYER M1 ;
		ANTENNAMAXAREACAR 16.533000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.010200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.151800 LAYER M2 ;
		ANTENNAMAXAREACAR 21.415000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.263800 LAYER M3 ;
		ANTENNAMAXAREACAR 316.698000 LAYER M3 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 141.896 17.375 141.976 ;
			LAYER M2 ;
			RECT 17.127 141.896 17.375 141.976 ;
			LAYER M3 ;
			RECT 17.127 141.896 17.375 141.976 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128800 LAYER M1 ;
		ANTENNAMAXAREACAR 16.533000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.010200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.151800 LAYER M2 ;
		ANTENNAMAXAREACAR 21.415000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.263800 LAYER M3 ;
		ANTENNAMAXAREACAR 316.698000 LAYER M3 ;
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.428 17.255 1.548 ;
			LAYER M4 ;
			RECT 0.120 1.932 17.255 2.052 ;
			LAYER M4 ;
			RECT 0.120 2.184 17.255 2.304 ;
			LAYER M4 ;
			RECT 0.120 3.444 17.255 3.564 ;
			LAYER M4 ;
			RECT 0.120 3.948 17.255 4.068 ;
			LAYER M4 ;
			RECT 0.120 4.200 17.255 4.320 ;
			LAYER M4 ;
			RECT 0.120 5.460 17.255 5.580 ;
			LAYER M4 ;
			RECT 0.120 5.964 17.255 6.084 ;
			LAYER M4 ;
			RECT 0.120 6.216 17.255 6.336 ;
			LAYER M4 ;
			RECT 0.120 7.476 17.255 7.596 ;
			LAYER M4 ;
			RECT 0.120 7.980 17.255 8.100 ;
			LAYER M4 ;
			RECT 0.120 8.232 17.255 8.352 ;
			LAYER M4 ;
			RECT 0.120 9.492 17.255 9.612 ;
			LAYER M4 ;
			RECT 0.120 9.996 17.255 10.116 ;
			LAYER M4 ;
			RECT 0.120 10.248 17.255 10.368 ;
			LAYER M4 ;
			RECT 0.120 11.508 17.255 11.628 ;
			LAYER M4 ;
			RECT 0.120 12.012 17.255 12.132 ;
			LAYER M4 ;
			RECT 0.120 12.264 17.255 12.384 ;
			LAYER M4 ;
			RECT 0.120 13.524 17.255 13.644 ;
			LAYER M4 ;
			RECT 0.120 14.028 17.255 14.148 ;
			LAYER M4 ;
			RECT 0.120 14.280 17.255 14.400 ;
			LAYER M4 ;
			RECT 0.120 15.540 17.255 15.660 ;
			LAYER M4 ;
			RECT 0.120 16.044 17.255 16.164 ;
			LAYER M4 ;
			RECT 0.120 16.296 17.255 16.416 ;
			LAYER M4 ;
			RECT 0.120 17.556 17.255 17.676 ;
			LAYER M4 ;
			RECT 0.120 18.060 17.255 18.180 ;
			LAYER M4 ;
			RECT 0.120 18.312 17.255 18.432 ;
			LAYER M4 ;
			RECT 0.120 19.572 17.255 19.692 ;
			LAYER M4 ;
			RECT 0.120 20.076 17.255 20.196 ;
			LAYER M4 ;
			RECT 0.120 20.328 17.255 20.448 ;
			LAYER M4 ;
			RECT 0.120 21.588 17.255 21.708 ;
			LAYER M4 ;
			RECT 0.120 22.092 17.255 22.212 ;
			LAYER M4 ;
			RECT 0.120 22.344 17.255 22.464 ;
			LAYER M4 ;
			RECT 0.120 23.604 17.255 23.724 ;
			LAYER M4 ;
			RECT 0.120 24.108 17.255 24.228 ;
			LAYER M4 ;
			RECT 0.120 24.360 17.255 24.480 ;
			LAYER M4 ;
			RECT 0.120 25.620 17.255 25.740 ;
			LAYER M4 ;
			RECT 0.120 26.124 17.255 26.244 ;
			LAYER M4 ;
			RECT 0.120 26.376 17.255 26.496 ;
			LAYER M4 ;
			RECT 0.120 27.636 17.255 27.756 ;
			LAYER M4 ;
			RECT 0.120 28.140 17.255 28.260 ;
			LAYER M4 ;
			RECT 0.120 28.392 17.255 28.512 ;
			LAYER M4 ;
			RECT 0.120 29.652 17.255 29.772 ;
			LAYER M4 ;
			RECT 0.120 30.156 17.255 30.276 ;
			LAYER M4 ;
			RECT 0.120 30.408 17.255 30.528 ;
			LAYER M4 ;
			RECT 0.120 31.668 17.255 31.788 ;
			LAYER M4 ;
			RECT 0.120 32.172 17.255 32.292 ;
			LAYER M4 ;
			RECT 0.120 32.424 17.255 32.544 ;
			LAYER M4 ;
			RECT 0.120 33.684 17.255 33.804 ;
			LAYER M4 ;
			RECT 0.120 34.188 17.255 34.308 ;
			LAYER M4 ;
			RECT 0.120 34.440 17.255 34.560 ;
			LAYER M4 ;
			RECT 0.120 35.700 17.255 35.820 ;
			LAYER M4 ;
			RECT 0.120 36.204 17.255 36.324 ;
			LAYER M4 ;
			RECT 0.120 36.456 17.255 36.576 ;
			LAYER M4 ;
			RECT 0.120 37.716 17.255 37.836 ;
			LAYER M4 ;
			RECT 0.120 38.220 17.255 38.340 ;
			LAYER M4 ;
			RECT 0.120 38.472 17.255 38.592 ;
			LAYER M4 ;
			RECT 0.120 39.732 17.255 39.852 ;
			LAYER M4 ;
			RECT 0.120 40.236 17.255 40.356 ;
			LAYER M4 ;
			RECT 0.120 40.488 17.255 40.608 ;
			LAYER M4 ;
			RECT 0.120 41.748 17.255 41.868 ;
			LAYER M4 ;
			RECT 0.120 42.252 17.255 42.372 ;
			LAYER M4 ;
			RECT 0.120 42.504 17.255 42.624 ;
			LAYER M4 ;
			RECT 0.120 43.764 17.255 43.884 ;
			LAYER M4 ;
			RECT 0.120 44.268 17.255 44.388 ;
			LAYER M4 ;
			RECT 0.120 44.520 17.255 44.640 ;
			LAYER M4 ;
			RECT 0.120 45.780 17.255 45.900 ;
			LAYER M4 ;
			RECT 0.120 46.284 17.255 46.404 ;
			LAYER M4 ;
			RECT 0.120 46.536 17.255 46.656 ;
			LAYER M4 ;
			RECT 0.120 47.796 17.255 47.916 ;
			LAYER M4 ;
			RECT 0.120 48.300 17.255 48.420 ;
			LAYER M4 ;
			RECT 0.120 48.552 17.255 48.672 ;
			LAYER M4 ;
			RECT 0.120 49.812 17.255 49.932 ;
			LAYER M4 ;
			RECT 0.120 50.316 17.255 50.436 ;
			LAYER M4 ;
			RECT 0.120 50.568 17.255 50.688 ;
			LAYER M4 ;
			RECT 0.120 51.828 17.255 51.948 ;
			LAYER M4 ;
			RECT 0.120 52.332 17.255 52.452 ;
			LAYER M4 ;
			RECT 0.120 52.584 17.255 52.704 ;
			LAYER M4 ;
			RECT 0.120 53.844 17.255 53.964 ;
			LAYER M4 ;
			RECT 0.120 54.348 17.255 54.468 ;
			LAYER M4 ;
			RECT 0.120 54.600 17.255 54.720 ;
			LAYER M4 ;
			RECT 0.120 55.860 17.255 55.980 ;
			LAYER M4 ;
			RECT 0.120 56.364 17.255 56.484 ;
			LAYER M4 ;
			RECT 0.120 56.616 17.255 56.736 ;
			LAYER M4 ;
			RECT 0.120 57.876 17.255 57.996 ;
			LAYER M4 ;
			RECT 0.120 58.380 17.255 58.500 ;
			LAYER M4 ;
			RECT 0.120 58.632 17.255 58.752 ;
			LAYER M4 ;
			RECT 0.120 59.892 17.255 60.012 ;
			LAYER M4 ;
			RECT 0.120 60.396 17.255 60.516 ;
			LAYER M4 ;
			RECT 0.120 60.648 17.255 60.768 ;
			LAYER M4 ;
			RECT 0.120 61.908 17.255 62.028 ;
			LAYER M4 ;
			RECT 0.120 62.412 17.255 62.532 ;
			LAYER M4 ;
			RECT 0.120 62.664 17.255 62.784 ;
			LAYER M4 ;
			RECT 0.120 63.924 17.255 64.044 ;
			LAYER M4 ;
			RECT 0.120 64.428 17.255 64.548 ;
			LAYER M4 ;
			RECT 0.120 64.680 17.255 64.800 ;
			LAYER M4 ;
			RECT 0.120 65.940 17.255 66.060 ;
			LAYER M4 ;
			RECT 0.120 66.444 17.255 66.564 ;
			LAYER M4 ;
			RECT 0.120 66.696 17.255 66.816 ;
			LAYER M4 ;
			RECT 0.120 67.956 17.255 68.076 ;
			LAYER M4 ;
			RECT 0.120 68.460 17.255 68.580 ;
			LAYER M4 ;
			RECT 0.120 68.712 17.255 68.832 ;
			LAYER M4 ;
			RECT 0.120 69.972 17.255 70.092 ;
			LAYER M4 ;
			RECT 0.120 70.476 17.255 70.596 ;
			LAYER M4 ;
			RECT 0.120 70.728 17.255 70.848 ;
			LAYER M4 ;
			RECT 0.120 71.988 17.255 72.108 ;
			LAYER M4 ;
			RECT 0.120 72.492 17.255 72.612 ;
			LAYER M4 ;
			RECT 0.120 72.744 17.255 72.864 ;
			LAYER M4 ;
			RECT 0.120 74.004 17.255 74.124 ;
			LAYER M4 ;
			RECT 0.120 74.508 17.255 74.628 ;
			LAYER M4 ;
			RECT 0.120 74.760 17.255 74.880 ;
			LAYER M4 ;
			RECT 0.120 76.020 17.255 76.140 ;
			LAYER M4 ;
			RECT 0.120 76.524 17.255 76.644 ;
			LAYER M4 ;
			RECT 0.120 76.776 17.255 76.896 ;
			LAYER M4 ;
			RECT 0.120 78.036 17.255 78.156 ;
			LAYER M4 ;
			RECT 0.120 78.540 17.255 78.660 ;
			LAYER M4 ;
			RECT 0.120 78.792 17.255 78.912 ;
			LAYER M4 ;
			RECT 0.120 80.052 17.255 80.172 ;
			LAYER M4 ;
			RECT 0.120 80.556 17.255 80.676 ;
			LAYER M4 ;
			RECT 0.120 80.808 17.255 80.928 ;
			LAYER M4 ;
			RECT 0.120 82.068 17.255 82.188 ;
			LAYER M4 ;
			RECT 0.120 82.572 17.255 82.692 ;
			LAYER M4 ;
			RECT 0.120 82.824 17.255 82.944 ;
			LAYER M4 ;
			RECT 0.120 84.084 17.255 84.204 ;
			LAYER M4 ;
			RECT 0.120 84.588 17.255 84.708 ;
			LAYER M4 ;
			RECT 0.120 84.840 17.255 84.960 ;
			LAYER M4 ;
			RECT 0.120 86.100 17.255 86.220 ;
			LAYER M4 ;
			RECT 0.120 86.604 17.255 86.724 ;
			LAYER M4 ;
			RECT 0.120 86.856 17.255 86.976 ;
			LAYER M4 ;
			RECT 0.120 88.116 17.255 88.236 ;
			LAYER M4 ;
			RECT 0.120 88.620 17.255 88.740 ;
			LAYER M4 ;
			RECT 0.120 88.872 17.255 88.992 ;
			LAYER M4 ;
			RECT 0.120 90.132 17.255 90.252 ;
			LAYER M4 ;
			RECT 0.120 90.636 17.255 90.756 ;
			LAYER M4 ;
			RECT 0.120 90.888 17.255 91.008 ;
			LAYER M4 ;
			RECT 0.120 92.148 17.255 92.268 ;
			LAYER M4 ;
			RECT 0.120 92.652 17.255 92.772 ;
			LAYER M4 ;
			RECT 0.120 92.904 17.255 93.024 ;
			LAYER M4 ;
			RECT 0.120 94.164 17.255 94.284 ;
			LAYER M4 ;
			RECT 0.120 94.668 17.255 94.788 ;
			LAYER M4 ;
			RECT 0.120 94.920 17.255 95.040 ;
			LAYER M4 ;
			RECT 0.120 96.180 17.255 96.300 ;
			LAYER M4 ;
			RECT 0.120 96.684 17.255 96.804 ;
			LAYER M4 ;
			RECT 0.120 96.936 17.255 97.056 ;
			LAYER M4 ;
			RECT 0.120 98.196 17.255 98.316 ;
			LAYER M4 ;
			RECT 0.120 98.700 17.255 98.820 ;
			LAYER M4 ;
			RECT 0.120 98.952 17.255 99.072 ;
			LAYER M4 ;
			RECT 0.120 100.212 17.255 100.332 ;
			LAYER M4 ;
			RECT 0.120 100.716 17.255 100.836 ;
			LAYER M4 ;
			RECT 0.120 100.968 17.255 101.088 ;
			LAYER M4 ;
			RECT 0.120 102.228 17.255 102.348 ;
			LAYER M4 ;
			RECT 0.120 102.732 17.255 102.852 ;
			LAYER M4 ;
			RECT 0.120 102.984 17.255 103.104 ;
			LAYER M4 ;
			RECT 0.120 104.244 17.255 104.364 ;
			LAYER M4 ;
			RECT 0.120 104.748 17.255 104.868 ;
			LAYER M4 ;
			RECT 0.120 105.000 17.255 105.120 ;
			LAYER M4 ;
			RECT 0.120 106.260 17.255 106.380 ;
			LAYER M4 ;
			RECT 0.120 106.764 17.255 106.884 ;
			LAYER M4 ;
			RECT 0.120 107.016 17.255 107.136 ;
			LAYER M4 ;
			RECT 0.120 108.276 17.255 108.396 ;
			LAYER M4 ;
			RECT 0.120 108.780 17.255 108.900 ;
			LAYER M4 ;
			RECT 0.120 109.032 17.255 109.152 ;
			LAYER M4 ;
			RECT 0.120 110.292 17.255 110.412 ;
			LAYER M4 ;
			RECT 0.120 110.796 17.255 110.916 ;
			LAYER M4 ;
			RECT 0.120 111.048 17.255 111.168 ;
			LAYER M4 ;
			RECT 0.120 112.308 17.255 112.428 ;
			LAYER M4 ;
			RECT 0.120 112.812 17.255 112.932 ;
			LAYER M4 ;
			RECT 0.120 113.064 17.255 113.184 ;
			LAYER M4 ;
			RECT 0.120 114.324 17.255 114.444 ;
			LAYER M4 ;
			RECT 0.120 114.828 17.255 114.948 ;
			LAYER M4 ;
			RECT 0.120 115.080 17.255 115.200 ;
			LAYER M4 ;
			RECT 0.120 116.340 17.255 116.460 ;
			LAYER M4 ;
			RECT 0.120 116.844 17.255 116.964 ;
			LAYER M4 ;
			RECT 0.120 117.096 17.255 117.216 ;
			LAYER M4 ;
			RECT 0.120 118.356 17.255 118.476 ;
			LAYER M4 ;
			RECT 0.120 118.860 17.255 118.980 ;
			LAYER M4 ;
			RECT 0.120 119.112 17.255 119.232 ;
			LAYER M4 ;
			RECT 0.120 120.372 17.255 120.492 ;
			LAYER M4 ;
			RECT 0.120 120.876 17.255 120.996 ;
			LAYER M4 ;
			RECT 0.120 121.128 17.255 121.248 ;
			LAYER M4 ;
			RECT 0.120 122.388 17.255 122.508 ;
			LAYER M4 ;
			RECT 0.120 122.892 17.255 123.012 ;
			LAYER M4 ;
			RECT 0.120 123.144 17.255 123.264 ;
			LAYER M4 ;
			RECT 0.120 124.404 17.255 124.524 ;
			LAYER M4 ;
			RECT 0.120 124.908 17.255 125.028 ;
			LAYER M4 ;
			RECT 0.120 125.160 17.255 125.280 ;
			LAYER M4 ;
			RECT 0.120 126.420 17.255 126.540 ;
			LAYER M4 ;
			RECT 0.120 126.924 17.255 127.044 ;
			LAYER M4 ;
			RECT 0.120 127.176 17.255 127.296 ;
			LAYER M4 ;
			RECT 0.120 128.436 17.255 128.556 ;
			LAYER M4 ;
			RECT 0.120 128.940 17.255 129.060 ;
			LAYER M4 ;
			RECT 0.120 129.192 17.255 129.312 ;
			LAYER M4 ;
			RECT 0.120 130.468 17.255 130.588 ;
			LAYER M4 ;
			RECT 0.120 131.092 17.255 131.212 ;
			LAYER M4 ;
			RECT 0.120 131.498 17.255 131.618 ;
			LAYER M4 ;
			RECT 0.120 131.958 17.255 132.078 ;
			LAYER M4 ;
			RECT 0.120 132.418 17.255 132.538 ;
			LAYER M4 ;
			RECT 0.120 132.878 17.255 132.998 ;
			LAYER M4 ;
			RECT 0.120 133.108 17.255 133.228 ;
			LAYER M4 ;
			RECT 0.120 133.500 17.255 133.620 ;
			LAYER M4 ;
			RECT 0.120 134.650 17.255 134.770 ;
			LAYER M4 ;
			RECT 0.120 135.332 17.255 135.452 ;
			LAYER M4 ;
			RECT 0.120 136.244 17.255 136.364 ;
			LAYER M4 ;
			RECT 0.120 137.423 17.255 137.543 ;
			LAYER M4 ;
			RECT 0.120 138.112 17.255 138.232 ;
			LAYER M4 ;
			RECT 0.120 138.572 17.255 138.692 ;
			LAYER M4 ;
			RECT 0.120 139.448 17.255 139.568 ;
			LAYER M4 ;
			RECT 0.120 139.908 17.255 140.028 ;
			LAYER M4 ;
			RECT 0.120 140.776 17.255 140.896 ;
			LAYER M4 ;
			RECT 0.120 141.210 17.255 141.330 ;
			LAYER M4 ;
			RECT 0.120 141.670 17.255 141.790 ;
			LAYER M4 ;
			RECT 0.120 142.080 17.255 142.200 ;
			LAYER M4 ;
			RECT 0.120 142.540 17.255 142.660 ;
			LAYER M4 ;
			RECT 0.120 143.316 17.255 143.436 ;
			LAYER M4 ;
			RECT 0.120 143.820 17.255 143.940 ;
			LAYER M4 ;
			RECT 0.120 144.072 17.255 144.192 ;
			LAYER M4 ;
			RECT 0.120 145.332 17.255 145.452 ;
			LAYER M4 ;
			RECT 0.120 145.836 17.255 145.956 ;
			LAYER M4 ;
			RECT 0.120 146.088 17.255 146.208 ;
			LAYER M4 ;
			RECT 0.120 147.348 17.255 147.468 ;
			LAYER M4 ;
			RECT 0.120 147.852 17.255 147.972 ;
			LAYER M4 ;
			RECT 0.120 148.104 17.255 148.224 ;
			LAYER M4 ;
			RECT 0.120 149.364 17.255 149.484 ;
			LAYER M4 ;
			RECT 0.120 149.868 17.255 149.988 ;
			LAYER M4 ;
			RECT 0.120 150.120 17.255 150.240 ;
			LAYER M4 ;
			RECT 0.120 151.380 17.255 151.500 ;
			LAYER M4 ;
			RECT 0.120 151.884 17.255 152.004 ;
			LAYER M4 ;
			RECT 0.120 152.136 17.255 152.256 ;
			LAYER M4 ;
			RECT 0.120 153.396 17.255 153.516 ;
			LAYER M4 ;
			RECT 0.120 153.900 17.255 154.020 ;
			LAYER M4 ;
			RECT 0.120 154.152 17.255 154.272 ;
			LAYER M4 ;
			RECT 0.120 155.412 17.255 155.532 ;
			LAYER M4 ;
			RECT 0.120 155.916 17.255 156.036 ;
			LAYER M4 ;
			RECT 0.120 156.168 17.255 156.288 ;
			LAYER M4 ;
			RECT 0.120 157.428 17.255 157.548 ;
			LAYER M4 ;
			RECT 0.120 157.932 17.255 158.052 ;
			LAYER M4 ;
			RECT 0.120 158.184 17.255 158.304 ;
			LAYER M4 ;
			RECT 0.120 159.444 17.255 159.564 ;
			LAYER M4 ;
			RECT 0.120 159.948 17.255 160.068 ;
			LAYER M4 ;
			RECT 0.120 160.200 17.255 160.320 ;
			LAYER M4 ;
			RECT 0.120 161.460 17.255 161.580 ;
			LAYER M4 ;
			RECT 0.120 161.964 17.255 162.084 ;
			LAYER M4 ;
			RECT 0.120 162.216 17.255 162.336 ;
			LAYER M4 ;
			RECT 0.120 163.476 17.255 163.596 ;
			LAYER M4 ;
			RECT 0.120 163.980 17.255 164.100 ;
			LAYER M4 ;
			RECT 0.120 164.232 17.255 164.352 ;
			LAYER M4 ;
			RECT 0.120 165.492 17.255 165.612 ;
			LAYER M4 ;
			RECT 0.120 165.996 17.255 166.116 ;
			LAYER M4 ;
			RECT 0.120 166.248 17.255 166.368 ;
			LAYER M4 ;
			RECT 0.120 167.508 17.255 167.628 ;
			LAYER M4 ;
			RECT 0.120 168.012 17.255 168.132 ;
			LAYER M4 ;
			RECT 0.120 168.264 17.255 168.384 ;
			LAYER M4 ;
			RECT 0.120 169.524 17.255 169.644 ;
			LAYER M4 ;
			RECT 0.120 170.028 17.255 170.148 ;
			LAYER M4 ;
			RECT 0.120 170.280 17.255 170.400 ;
			LAYER M4 ;
			RECT 0.120 171.540 17.255 171.660 ;
			LAYER M4 ;
			RECT 0.120 172.044 17.255 172.164 ;
			LAYER M4 ;
			RECT 0.120 172.296 17.255 172.416 ;
			LAYER M4 ;
			RECT 0.120 173.556 17.255 173.676 ;
			LAYER M4 ;
			RECT 0.120 174.060 17.255 174.180 ;
			LAYER M4 ;
			RECT 0.120 174.312 17.255 174.432 ;
			LAYER M4 ;
			RECT 0.120 175.572 17.255 175.692 ;
			LAYER M4 ;
			RECT 0.120 176.076 17.255 176.196 ;
			LAYER M4 ;
			RECT 0.120 176.328 17.255 176.448 ;
			LAYER M4 ;
			RECT 0.120 177.588 17.255 177.708 ;
			LAYER M4 ;
			RECT 0.120 178.092 17.255 178.212 ;
			LAYER M4 ;
			RECT 0.120 178.344 17.255 178.464 ;
			LAYER M4 ;
			RECT 0.120 179.604 17.255 179.724 ;
			LAYER M4 ;
			RECT 0.120 180.108 17.255 180.228 ;
			LAYER M4 ;
			RECT 0.120 180.360 17.255 180.480 ;
			LAYER M4 ;
			RECT 0.120 181.620 17.255 181.740 ;
			LAYER M4 ;
			RECT 0.120 182.124 17.255 182.244 ;
			LAYER M4 ;
			RECT 0.120 182.376 17.255 182.496 ;
			LAYER M4 ;
			RECT 0.120 183.636 17.255 183.756 ;
			LAYER M4 ;
			RECT 0.120 184.140 17.255 184.260 ;
			LAYER M4 ;
			RECT 0.120 184.392 17.255 184.512 ;
			LAYER M4 ;
			RECT 0.120 185.652 17.255 185.772 ;
			LAYER M4 ;
			RECT 0.120 186.156 17.255 186.276 ;
			LAYER M4 ;
			RECT 0.120 186.408 17.255 186.528 ;
			LAYER M4 ;
			RECT 0.120 187.668 17.255 187.788 ;
			LAYER M4 ;
			RECT 0.120 188.172 17.255 188.292 ;
			LAYER M4 ;
			RECT 0.120 188.424 17.255 188.544 ;
			LAYER M4 ;
			RECT 0.120 189.684 17.255 189.804 ;
			LAYER M4 ;
			RECT 0.120 190.188 17.255 190.308 ;
			LAYER M4 ;
			RECT 0.120 190.440 17.255 190.560 ;
			LAYER M4 ;
			RECT 0.120 191.700 17.255 191.820 ;
			LAYER M4 ;
			RECT 0.120 192.204 17.255 192.324 ;
			LAYER M4 ;
			RECT 0.120 192.456 17.255 192.576 ;
			LAYER M4 ;
			RECT 0.120 193.716 17.255 193.836 ;
			LAYER M4 ;
			RECT 0.120 194.220 17.255 194.340 ;
			LAYER M4 ;
			RECT 0.120 194.472 17.255 194.592 ;
			LAYER M4 ;
			RECT 0.120 195.732 17.255 195.852 ;
			LAYER M4 ;
			RECT 0.120 196.236 17.255 196.356 ;
			LAYER M4 ;
			RECT 0.120 196.488 17.255 196.608 ;
			LAYER M4 ;
			RECT 0.120 197.748 17.255 197.868 ;
			LAYER M4 ;
			RECT 0.120 198.252 17.255 198.372 ;
			LAYER M4 ;
			RECT 0.120 198.504 17.255 198.624 ;
			LAYER M4 ;
			RECT 0.120 199.764 17.255 199.884 ;
			LAYER M4 ;
			RECT 0.120 200.268 17.255 200.388 ;
			LAYER M4 ;
			RECT 0.120 200.520 17.255 200.640 ;
			LAYER M4 ;
			RECT 0.120 201.780 17.255 201.900 ;
			LAYER M4 ;
			RECT 0.120 202.284 17.255 202.404 ;
			LAYER M4 ;
			RECT 0.120 202.536 17.255 202.656 ;
			LAYER M4 ;
			RECT 0.120 203.796 17.255 203.916 ;
			LAYER M4 ;
			RECT 0.120 204.300 17.255 204.420 ;
			LAYER M4 ;
			RECT 0.120 204.552 17.255 204.672 ;
			LAYER M4 ;
			RECT 0.120 205.812 17.255 205.932 ;
			LAYER M4 ;
			RECT 0.120 206.316 17.255 206.436 ;
			LAYER M4 ;
			RECT 0.120 206.568 17.255 206.688 ;
			LAYER M4 ;
			RECT 0.120 207.828 17.255 207.948 ;
			LAYER M4 ;
			RECT 0.120 208.332 17.255 208.452 ;
			LAYER M4 ;
			RECT 0.120 208.584 17.255 208.704 ;
			LAYER M4 ;
			RECT 0.120 209.844 17.255 209.964 ;
			LAYER M4 ;
			RECT 0.120 210.348 17.255 210.468 ;
			LAYER M4 ;
			RECT 0.120 210.600 17.255 210.720 ;
			LAYER M4 ;
			RECT 0.120 211.860 17.255 211.980 ;
			LAYER M4 ;
			RECT 0.120 212.364 17.255 212.484 ;
			LAYER M4 ;
			RECT 0.120 212.616 17.255 212.736 ;
			LAYER M4 ;
			RECT 0.120 213.876 17.255 213.996 ;
			LAYER M4 ;
			RECT 0.120 214.380 17.255 214.500 ;
			LAYER M4 ;
			RECT 0.120 214.632 17.255 214.752 ;
			LAYER M4 ;
			RECT 0.120 215.892 17.255 216.012 ;
			LAYER M4 ;
			RECT 0.120 216.396 17.255 216.516 ;
			LAYER M4 ;
			RECT 0.120 216.648 17.255 216.768 ;
			LAYER M4 ;
			RECT 0.120 217.908 17.255 218.028 ;
			LAYER M4 ;
			RECT 0.120 218.412 17.255 218.532 ;
			LAYER M4 ;
			RECT 0.120 218.664 17.255 218.784 ;
			LAYER M4 ;
			RECT 0.120 219.924 17.255 220.044 ;
			LAYER M4 ;
			RECT 0.120 220.428 17.255 220.548 ;
			LAYER M4 ;
			RECT 0.120 220.680 17.255 220.800 ;
			LAYER M4 ;
			RECT 0.120 221.940 17.255 222.060 ;
			LAYER M4 ;
			RECT 0.120 222.444 17.255 222.564 ;
			LAYER M4 ;
			RECT 0.120 222.696 17.255 222.816 ;
			LAYER M4 ;
			RECT 0.120 223.956 17.255 224.076 ;
			LAYER M4 ;
			RECT 0.120 224.460 17.255 224.580 ;
			LAYER M4 ;
			RECT 0.120 224.712 17.255 224.832 ;
			LAYER M4 ;
			RECT 0.120 225.972 17.255 226.092 ;
			LAYER M4 ;
			RECT 0.120 226.476 17.255 226.596 ;
			LAYER M4 ;
			RECT 0.120 226.728 17.255 226.848 ;
			LAYER M4 ;
			RECT 0.120 227.988 17.255 228.108 ;
			LAYER M4 ;
			RECT 0.120 228.492 17.255 228.612 ;
			LAYER M4 ;
			RECT 0.120 228.744 17.255 228.864 ;
			LAYER M4 ;
			RECT 0.120 230.004 17.255 230.124 ;
			LAYER M4 ;
			RECT 0.120 230.508 17.255 230.628 ;
			LAYER M4 ;
			RECT 0.120 230.760 17.255 230.880 ;
			LAYER M4 ;
			RECT 0.120 232.020 17.255 232.140 ;
			LAYER M4 ;
			RECT 0.120 232.524 17.255 232.644 ;
			LAYER M4 ;
			RECT 0.120 232.776 17.255 232.896 ;
			LAYER M4 ;
			RECT 0.120 234.036 17.255 234.156 ;
			LAYER M4 ;
			RECT 0.120 234.540 17.255 234.660 ;
			LAYER M4 ;
			RECT 0.120 234.792 17.255 234.912 ;
			LAYER M4 ;
			RECT 0.120 236.052 17.255 236.172 ;
			LAYER M4 ;
			RECT 0.120 236.556 17.255 236.676 ;
			LAYER M4 ;
			RECT 0.120 236.808 17.255 236.928 ;
			LAYER M4 ;
			RECT 0.120 238.068 17.255 238.188 ;
			LAYER M4 ;
			RECT 0.120 238.572 17.255 238.692 ;
			LAYER M4 ;
			RECT 0.120 238.824 17.255 238.944 ;
			LAYER M4 ;
			RECT 0.120 240.084 17.255 240.204 ;
			LAYER M4 ;
			RECT 0.120 240.588 17.255 240.708 ;
			LAYER M4 ;
			RECT 0.120 240.840 17.255 240.960 ;
			LAYER M4 ;
			RECT 0.120 242.100 17.255 242.220 ;
			LAYER M4 ;
			RECT 0.120 242.604 17.255 242.724 ;
			LAYER M4 ;
			RECT 0.120 242.856 17.255 242.976 ;
			LAYER M4 ;
			RECT 0.120 244.116 17.255 244.236 ;
			LAYER M4 ;
			RECT 0.120 244.620 17.255 244.740 ;
			LAYER M4 ;
			RECT 0.120 244.872 17.255 244.992 ;
			LAYER M4 ;
			RECT 0.120 246.132 17.255 246.252 ;
			LAYER M4 ;
			RECT 0.120 246.636 17.255 246.756 ;
			LAYER M4 ;
			RECT 0.120 246.888 17.255 247.008 ;
			LAYER M4 ;
			RECT 0.120 248.148 17.255 248.268 ;
			LAYER M4 ;
			RECT 0.120 248.652 17.255 248.772 ;
			LAYER M4 ;
			RECT 0.120 248.904 17.255 249.024 ;
			LAYER M4 ;
			RECT 0.120 250.164 17.255 250.284 ;
			LAYER M4 ;
			RECT 0.120 250.668 17.255 250.788 ;
			LAYER M4 ;
			RECT 0.120 250.920 17.255 251.040 ;
			LAYER M4 ;
			RECT 0.120 252.180 17.255 252.300 ;
			LAYER M4 ;
			RECT 0.120 252.684 17.255 252.804 ;
			LAYER M4 ;
			RECT 0.120 252.936 17.255 253.056 ;
			LAYER M4 ;
			RECT 0.120 254.196 17.255 254.316 ;
			LAYER M4 ;
			RECT 0.120 254.700 17.255 254.820 ;
			LAYER M4 ;
			RECT 0.120 254.952 17.255 255.072 ;
			LAYER M4 ;
			RECT 0.120 256.212 17.255 256.332 ;
			LAYER M4 ;
			RECT 0.120 256.716 17.255 256.836 ;
			LAYER M4 ;
			RECT 0.120 256.968 17.255 257.088 ;
			LAYER M4 ;
			RECT 0.120 258.228 17.255 258.348 ;
			LAYER M4 ;
			RECT 0.120 258.732 17.255 258.852 ;
			LAYER M4 ;
			RECT 0.120 258.984 17.255 259.104 ;
			LAYER M4 ;
			RECT 0.120 260.244 17.255 260.364 ;
			LAYER M4 ;
			RECT 0.120 260.748 17.255 260.868 ;
			LAYER M4 ;
			RECT 0.120 261.000 17.255 261.120 ;
			LAYER M4 ;
			RECT 0.120 262.260 17.255 262.380 ;
			LAYER M4 ;
			RECT 0.120 262.764 17.255 262.884 ;
			LAYER M4 ;
			RECT 0.120 263.016 17.255 263.136 ;
			LAYER M4 ;
			RECT 0.120 264.276 17.255 264.396 ;
			LAYER M4 ;
			RECT 0.120 264.780 17.255 264.900 ;
			LAYER M4 ;
			RECT 0.120 265.032 17.255 265.152 ;
			LAYER M4 ;
			RECT 0.120 266.292 17.255 266.412 ;
			LAYER M4 ;
			RECT 0.120 266.796 17.255 266.916 ;
			LAYER M4 ;
			RECT 0.120 267.048 17.255 267.168 ;
			LAYER M4 ;
			RECT 0.120 268.308 17.255 268.428 ;
			LAYER M4 ;
			RECT 0.120 268.812 17.255 268.932 ;
			LAYER M4 ;
			RECT 0.120 269.064 17.255 269.184 ;
			LAYER M4 ;
			RECT 0.120 270.324 17.255 270.444 ;
			LAYER M4 ;
			RECT 0.120 270.828 17.255 270.948 ;
			LAYER M4 ;
			RECT 0.120 271.080 17.255 271.200 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.176 17.255 1.296 ;
			LAYER M4 ;
			RECT 0.120 1.680 17.255 1.800 ;
			LAYER M4 ;
			RECT 0.120 2.688 17.255 2.808 ;
			LAYER M4 ;
			RECT 0.120 3.192 17.255 3.312 ;
			LAYER M4 ;
			RECT 0.120 3.696 17.255 3.816 ;
			LAYER M4 ;
			RECT 0.120 4.704 17.255 4.824 ;
			LAYER M4 ;
			RECT 0.120 5.208 17.255 5.328 ;
			LAYER M4 ;
			RECT 0.120 5.712 17.255 5.832 ;
			LAYER M4 ;
			RECT 0.120 6.720 17.255 6.840 ;
			LAYER M4 ;
			RECT 0.120 7.224 17.255 7.344 ;
			LAYER M4 ;
			RECT 0.120 7.728 17.255 7.848 ;
			LAYER M4 ;
			RECT 0.120 8.736 17.255 8.856 ;
			LAYER M4 ;
			RECT 0.120 9.240 17.255 9.360 ;
			LAYER M4 ;
			RECT 0.120 9.744 17.255 9.864 ;
			LAYER M4 ;
			RECT 0.120 10.752 17.255 10.872 ;
			LAYER M4 ;
			RECT 0.120 11.256 17.255 11.376 ;
			LAYER M4 ;
			RECT 0.120 11.760 17.255 11.880 ;
			LAYER M4 ;
			RECT 0.120 12.768 17.255 12.888 ;
			LAYER M4 ;
			RECT 0.120 13.272 17.255 13.392 ;
			LAYER M4 ;
			RECT 0.120 13.776 17.255 13.896 ;
			LAYER M4 ;
			RECT 0.120 14.784 17.255 14.904 ;
			LAYER M4 ;
			RECT 0.120 15.288 17.255 15.408 ;
			LAYER M4 ;
			RECT 0.120 15.792 17.255 15.912 ;
			LAYER M4 ;
			RECT 0.120 16.800 17.255 16.920 ;
			LAYER M4 ;
			RECT 0.120 17.304 17.255 17.424 ;
			LAYER M4 ;
			RECT 0.120 17.808 17.255 17.928 ;
			LAYER M4 ;
			RECT 0.120 18.816 17.255 18.936 ;
			LAYER M4 ;
			RECT 0.120 19.320 17.255 19.440 ;
			LAYER M4 ;
			RECT 0.120 19.824 17.255 19.944 ;
			LAYER M4 ;
			RECT 0.120 20.832 17.255 20.952 ;
			LAYER M4 ;
			RECT 0.120 21.336 17.255 21.456 ;
			LAYER M4 ;
			RECT 0.120 21.840 17.255 21.960 ;
			LAYER M4 ;
			RECT 0.120 22.848 17.255 22.968 ;
			LAYER M4 ;
			RECT 0.120 23.352 17.255 23.472 ;
			LAYER M4 ;
			RECT 0.120 23.856 17.255 23.976 ;
			LAYER M4 ;
			RECT 0.120 24.864 17.255 24.984 ;
			LAYER M4 ;
			RECT 0.120 25.368 17.255 25.488 ;
			LAYER M4 ;
			RECT 0.120 25.872 17.255 25.992 ;
			LAYER M4 ;
			RECT 0.120 26.880 17.255 27.000 ;
			LAYER M4 ;
			RECT 0.120 27.384 17.255 27.504 ;
			LAYER M4 ;
			RECT 0.120 27.888 17.255 28.008 ;
			LAYER M4 ;
			RECT 0.120 28.896 17.255 29.016 ;
			LAYER M4 ;
			RECT 0.120 29.400 17.255 29.520 ;
			LAYER M4 ;
			RECT 0.120 29.904 17.255 30.024 ;
			LAYER M4 ;
			RECT 0.120 30.912 17.255 31.032 ;
			LAYER M4 ;
			RECT 0.120 31.416 17.255 31.536 ;
			LAYER M4 ;
			RECT 0.120 31.920 17.255 32.040 ;
			LAYER M4 ;
			RECT 0.120 32.928 17.255 33.048 ;
			LAYER M4 ;
			RECT 0.120 33.432 17.255 33.552 ;
			LAYER M4 ;
			RECT 0.120 33.936 17.255 34.056 ;
			LAYER M4 ;
			RECT 0.120 34.944 17.255 35.064 ;
			LAYER M4 ;
			RECT 0.120 35.448 17.255 35.568 ;
			LAYER M4 ;
			RECT 0.120 35.952 17.255 36.072 ;
			LAYER M4 ;
			RECT 0.120 36.960 17.255 37.080 ;
			LAYER M4 ;
			RECT 0.120 37.464 17.255 37.584 ;
			LAYER M4 ;
			RECT 0.120 37.968 17.255 38.088 ;
			LAYER M4 ;
			RECT 0.120 38.976 17.255 39.096 ;
			LAYER M4 ;
			RECT 0.120 39.480 17.255 39.600 ;
			LAYER M4 ;
			RECT 0.120 39.984 17.255 40.104 ;
			LAYER M4 ;
			RECT 0.120 40.992 17.255 41.112 ;
			LAYER M4 ;
			RECT 0.120 41.496 17.255 41.616 ;
			LAYER M4 ;
			RECT 0.120 42.000 17.255 42.120 ;
			LAYER M4 ;
			RECT 0.120 43.008 17.255 43.128 ;
			LAYER M4 ;
			RECT 0.120 43.512 17.255 43.632 ;
			LAYER M4 ;
			RECT 0.120 44.016 17.255 44.136 ;
			LAYER M4 ;
			RECT 0.120 45.024 17.255 45.144 ;
			LAYER M4 ;
			RECT 0.120 45.528 17.255 45.648 ;
			LAYER M4 ;
			RECT 0.120 46.032 17.255 46.152 ;
			LAYER M4 ;
			RECT 0.120 47.040 17.255 47.160 ;
			LAYER M4 ;
			RECT 0.120 47.544 17.255 47.664 ;
			LAYER M4 ;
			RECT 0.120 48.048 17.255 48.168 ;
			LAYER M4 ;
			RECT 0.120 49.056 17.255 49.176 ;
			LAYER M4 ;
			RECT 0.120 49.560 17.255 49.680 ;
			LAYER M4 ;
			RECT 0.120 50.064 17.255 50.184 ;
			LAYER M4 ;
			RECT 0.120 51.072 17.255 51.192 ;
			LAYER M4 ;
			RECT 0.120 51.576 17.255 51.696 ;
			LAYER M4 ;
			RECT 0.120 52.080 17.255 52.200 ;
			LAYER M4 ;
			RECT 0.120 53.088 17.255 53.208 ;
			LAYER M4 ;
			RECT 0.120 53.592 17.255 53.712 ;
			LAYER M4 ;
			RECT 0.120 54.096 17.255 54.216 ;
			LAYER M4 ;
			RECT 0.120 55.104 17.255 55.224 ;
			LAYER M4 ;
			RECT 0.120 55.608 17.255 55.728 ;
			LAYER M4 ;
			RECT 0.120 56.112 17.255 56.232 ;
			LAYER M4 ;
			RECT 0.120 57.120 17.255 57.240 ;
			LAYER M4 ;
			RECT 0.120 57.624 17.255 57.744 ;
			LAYER M4 ;
			RECT 0.120 58.128 17.255 58.248 ;
			LAYER M4 ;
			RECT 0.120 59.136 17.255 59.256 ;
			LAYER M4 ;
			RECT 0.120 59.640 17.255 59.760 ;
			LAYER M4 ;
			RECT 0.120 60.144 17.255 60.264 ;
			LAYER M4 ;
			RECT 0.120 61.152 17.255 61.272 ;
			LAYER M4 ;
			RECT 0.120 61.656 17.255 61.776 ;
			LAYER M4 ;
			RECT 0.120 62.160 17.255 62.280 ;
			LAYER M4 ;
			RECT 0.120 63.168 17.255 63.288 ;
			LAYER M4 ;
			RECT 0.120 63.672 17.255 63.792 ;
			LAYER M4 ;
			RECT 0.120 64.176 17.255 64.296 ;
			LAYER M4 ;
			RECT 0.120 65.184 17.255 65.304 ;
			LAYER M4 ;
			RECT 0.120 65.688 17.255 65.808 ;
			LAYER M4 ;
			RECT 0.120 66.192 17.255 66.312 ;
			LAYER M4 ;
			RECT 0.120 67.200 17.255 67.320 ;
			LAYER M4 ;
			RECT 0.120 67.704 17.255 67.824 ;
			LAYER M4 ;
			RECT 0.120 68.208 17.255 68.328 ;
			LAYER M4 ;
			RECT 0.120 69.216 17.255 69.336 ;
			LAYER M4 ;
			RECT 0.120 69.720 17.255 69.840 ;
			LAYER M4 ;
			RECT 0.120 70.224 17.255 70.344 ;
			LAYER M4 ;
			RECT 0.120 71.232 17.255 71.352 ;
			LAYER M4 ;
			RECT 0.120 71.736 17.255 71.856 ;
			LAYER M4 ;
			RECT 0.120 72.240 17.255 72.360 ;
			LAYER M4 ;
			RECT 0.120 73.248 17.255 73.368 ;
			LAYER M4 ;
			RECT 0.120 73.752 17.255 73.872 ;
			LAYER M4 ;
			RECT 0.120 74.256 17.255 74.376 ;
			LAYER M4 ;
			RECT 0.120 75.264 17.255 75.384 ;
			LAYER M4 ;
			RECT 0.120 75.768 17.255 75.888 ;
			LAYER M4 ;
			RECT 0.120 76.272 17.255 76.392 ;
			LAYER M4 ;
			RECT 0.120 77.280 17.255 77.400 ;
			LAYER M4 ;
			RECT 0.120 77.784 17.255 77.904 ;
			LAYER M4 ;
			RECT 0.120 78.288 17.255 78.408 ;
			LAYER M4 ;
			RECT 0.120 79.296 17.255 79.416 ;
			LAYER M4 ;
			RECT 0.120 79.800 17.255 79.920 ;
			LAYER M4 ;
			RECT 0.120 80.304 17.255 80.424 ;
			LAYER M4 ;
			RECT 0.120 81.312 17.255 81.432 ;
			LAYER M4 ;
			RECT 0.120 81.816 17.255 81.936 ;
			LAYER M4 ;
			RECT 0.120 82.320 17.255 82.440 ;
			LAYER M4 ;
			RECT 0.120 83.328 17.255 83.448 ;
			LAYER M4 ;
			RECT 0.120 83.832 17.255 83.952 ;
			LAYER M4 ;
			RECT 0.120 84.336 17.255 84.456 ;
			LAYER M4 ;
			RECT 0.120 85.344 17.255 85.464 ;
			LAYER M4 ;
			RECT 0.120 85.848 17.255 85.968 ;
			LAYER M4 ;
			RECT 0.120 86.352 17.255 86.472 ;
			LAYER M4 ;
			RECT 0.120 87.360 17.255 87.480 ;
			LAYER M4 ;
			RECT 0.120 87.864 17.255 87.984 ;
			LAYER M4 ;
			RECT 0.120 88.368 17.255 88.488 ;
			LAYER M4 ;
			RECT 0.120 89.376 17.255 89.496 ;
			LAYER M4 ;
			RECT 0.120 89.880 17.255 90.000 ;
			LAYER M4 ;
			RECT 0.120 90.384 17.255 90.504 ;
			LAYER M4 ;
			RECT 0.120 91.392 17.255 91.512 ;
			LAYER M4 ;
			RECT 0.120 91.896 17.255 92.016 ;
			LAYER M4 ;
			RECT 0.120 92.400 17.255 92.520 ;
			LAYER M4 ;
			RECT 0.120 93.408 17.255 93.528 ;
			LAYER M4 ;
			RECT 0.120 93.912 17.255 94.032 ;
			LAYER M4 ;
			RECT 0.120 94.416 17.255 94.536 ;
			LAYER M4 ;
			RECT 0.120 95.424 17.255 95.544 ;
			LAYER M4 ;
			RECT 0.120 95.928 17.255 96.048 ;
			LAYER M4 ;
			RECT 0.120 96.432 17.255 96.552 ;
			LAYER M4 ;
			RECT 0.120 97.440 17.255 97.560 ;
			LAYER M4 ;
			RECT 0.120 97.944 17.255 98.064 ;
			LAYER M4 ;
			RECT 0.120 98.448 17.255 98.568 ;
			LAYER M4 ;
			RECT 0.120 99.456 17.255 99.576 ;
			LAYER M4 ;
			RECT 0.120 99.960 17.255 100.080 ;
			LAYER M4 ;
			RECT 0.120 100.464 17.255 100.584 ;
			LAYER M4 ;
			RECT 0.120 101.472 17.255 101.592 ;
			LAYER M4 ;
			RECT 0.120 101.976 17.255 102.096 ;
			LAYER M4 ;
			RECT 0.120 102.480 17.255 102.600 ;
			LAYER M4 ;
			RECT 0.120 103.488 17.255 103.608 ;
			LAYER M4 ;
			RECT 0.120 103.992 17.255 104.112 ;
			LAYER M4 ;
			RECT 0.120 104.496 17.255 104.616 ;
			LAYER M4 ;
			RECT 0.120 105.504 17.255 105.624 ;
			LAYER M4 ;
			RECT 0.120 106.008 17.255 106.128 ;
			LAYER M4 ;
			RECT 0.120 106.512 17.255 106.632 ;
			LAYER M4 ;
			RECT 0.120 107.520 17.255 107.640 ;
			LAYER M4 ;
			RECT 0.120 108.024 17.255 108.144 ;
			LAYER M4 ;
			RECT 0.120 108.528 17.255 108.648 ;
			LAYER M4 ;
			RECT 0.120 109.536 17.255 109.656 ;
			LAYER M4 ;
			RECT 0.120 110.040 17.255 110.160 ;
			LAYER M4 ;
			RECT 0.120 110.544 17.255 110.664 ;
			LAYER M4 ;
			RECT 0.120 111.552 17.255 111.672 ;
			LAYER M4 ;
			RECT 0.120 112.056 17.255 112.176 ;
			LAYER M4 ;
			RECT 0.120 112.560 17.255 112.680 ;
			LAYER M4 ;
			RECT 0.120 113.568 17.255 113.688 ;
			LAYER M4 ;
			RECT 0.120 114.072 17.255 114.192 ;
			LAYER M4 ;
			RECT 0.120 114.576 17.255 114.696 ;
			LAYER M4 ;
			RECT 0.120 115.584 17.255 115.704 ;
			LAYER M4 ;
			RECT 0.120 116.088 17.255 116.208 ;
			LAYER M4 ;
			RECT 0.120 116.592 17.255 116.712 ;
			LAYER M4 ;
			RECT 0.120 117.600 17.255 117.720 ;
			LAYER M4 ;
			RECT 0.120 118.104 17.255 118.224 ;
			LAYER M4 ;
			RECT 0.120 118.608 17.255 118.728 ;
			LAYER M4 ;
			RECT 0.120 119.616 17.255 119.736 ;
			LAYER M4 ;
			RECT 0.120 120.120 17.255 120.240 ;
			LAYER M4 ;
			RECT 0.120 120.624 17.255 120.744 ;
			LAYER M4 ;
			RECT 0.120 121.632 17.255 121.752 ;
			LAYER M4 ;
			RECT 0.120 122.136 17.255 122.256 ;
			LAYER M4 ;
			RECT 0.120 122.640 17.255 122.760 ;
			LAYER M4 ;
			RECT 0.120 123.648 17.255 123.768 ;
			LAYER M4 ;
			RECT 0.120 124.152 17.255 124.272 ;
			LAYER M4 ;
			RECT 0.120 124.656 17.255 124.776 ;
			LAYER M4 ;
			RECT 0.120 125.664 17.255 125.784 ;
			LAYER M4 ;
			RECT 0.120 126.168 17.255 126.288 ;
			LAYER M4 ;
			RECT 0.120 126.672 17.255 126.792 ;
			LAYER M4 ;
			RECT 0.120 127.680 17.255 127.800 ;
			LAYER M4 ;
			RECT 0.120 128.184 17.255 128.304 ;
			LAYER M4 ;
			RECT 0.120 128.688 17.255 128.808 ;
			LAYER M4 ;
			RECT 0.120 129.696 17.255 129.816 ;
			LAYER M4 ;
			RECT 0.120 130.862 17.255 130.982 ;
			LAYER M4 ;
			RECT 0.120 131.728 17.255 131.848 ;
			LAYER M4 ;
			RECT 0.120 132.188 17.255 132.308 ;
			LAYER M4 ;
			RECT 0.120 132.648 17.255 132.768 ;
			LAYER M4 ;
			RECT 0.120 133.730 17.255 133.850 ;
			LAYER M4 ;
			RECT 0.120 134.420 17.255 134.540 ;
			LAYER M4 ;
			RECT 0.120 135.562 17.255 135.682 ;
			LAYER M4 ;
			RECT 0.120 136.474 17.255 136.594 ;
			LAYER M4 ;
			RECT 0.120 137.193 17.255 137.313 ;
			LAYER M4 ;
			RECT 0.120 138.342 17.255 138.462 ;
			LAYER M4 ;
			RECT 0.120 138.802 17.255 138.922 ;
			LAYER M4 ;
			RECT 0.120 139.218 17.255 139.338 ;
			LAYER M4 ;
			RECT 0.120 139.678 17.255 139.798 ;
			LAYER M4 ;
			RECT 0.120 140.138 17.255 140.258 ;
			LAYER M4 ;
			RECT 0.120 140.546 17.255 140.666 ;
			LAYER M4 ;
			RECT 0.120 141.440 17.255 141.560 ;
			LAYER M4 ;
			RECT 0.120 142.310 17.255 142.430 ;
			LAYER M4 ;
			RECT 0.120 143.064 17.255 143.184 ;
			LAYER M4 ;
			RECT 0.120 143.568 17.255 143.688 ;
			LAYER M4 ;
			RECT 0.120 144.576 17.255 144.696 ;
			LAYER M4 ;
			RECT 0.120 145.080 17.255 145.200 ;
			LAYER M4 ;
			RECT 0.120 145.584 17.255 145.704 ;
			LAYER M4 ;
			RECT 0.120 146.592 17.255 146.712 ;
			LAYER M4 ;
			RECT 0.120 147.096 17.255 147.216 ;
			LAYER M4 ;
			RECT 0.120 147.600 17.255 147.720 ;
			LAYER M4 ;
			RECT 0.120 148.608 17.255 148.728 ;
			LAYER M4 ;
			RECT 0.120 149.112 17.255 149.232 ;
			LAYER M4 ;
			RECT 0.120 149.616 17.255 149.736 ;
			LAYER M4 ;
			RECT 0.120 150.624 17.255 150.744 ;
			LAYER M4 ;
			RECT 0.120 151.128 17.255 151.248 ;
			LAYER M4 ;
			RECT 0.120 151.632 17.255 151.752 ;
			LAYER M4 ;
			RECT 0.120 152.640 17.255 152.760 ;
			LAYER M4 ;
			RECT 0.120 153.144 17.255 153.264 ;
			LAYER M4 ;
			RECT 0.120 153.648 17.255 153.768 ;
			LAYER M4 ;
			RECT 0.120 154.656 17.255 154.776 ;
			LAYER M4 ;
			RECT 0.120 155.160 17.255 155.280 ;
			LAYER M4 ;
			RECT 0.120 155.664 17.255 155.784 ;
			LAYER M4 ;
			RECT 0.120 156.672 17.255 156.792 ;
			LAYER M4 ;
			RECT 0.120 157.176 17.255 157.296 ;
			LAYER M4 ;
			RECT 0.120 157.680 17.255 157.800 ;
			LAYER M4 ;
			RECT 0.120 158.688 17.255 158.808 ;
			LAYER M4 ;
			RECT 0.120 159.192 17.255 159.312 ;
			LAYER M4 ;
			RECT 0.120 159.696 17.255 159.816 ;
			LAYER M4 ;
			RECT 0.120 160.704 17.255 160.824 ;
			LAYER M4 ;
			RECT 0.120 161.208 17.255 161.328 ;
			LAYER M4 ;
			RECT 0.120 161.712 17.255 161.832 ;
			LAYER M4 ;
			RECT 0.120 162.720 17.255 162.840 ;
			LAYER M4 ;
			RECT 0.120 163.224 17.255 163.344 ;
			LAYER M4 ;
			RECT 0.120 163.728 17.255 163.848 ;
			LAYER M4 ;
			RECT 0.120 164.736 17.255 164.856 ;
			LAYER M4 ;
			RECT 0.120 165.240 17.255 165.360 ;
			LAYER M4 ;
			RECT 0.120 165.744 17.255 165.864 ;
			LAYER M4 ;
			RECT 0.120 166.752 17.255 166.872 ;
			LAYER M4 ;
			RECT 0.120 167.256 17.255 167.376 ;
			LAYER M4 ;
			RECT 0.120 167.760 17.255 167.880 ;
			LAYER M4 ;
			RECT 0.120 168.768 17.255 168.888 ;
			LAYER M4 ;
			RECT 0.120 169.272 17.255 169.392 ;
			LAYER M4 ;
			RECT 0.120 169.776 17.255 169.896 ;
			LAYER M4 ;
			RECT 0.120 170.784 17.255 170.904 ;
			LAYER M4 ;
			RECT 0.120 171.288 17.255 171.408 ;
			LAYER M4 ;
			RECT 0.120 171.792 17.255 171.912 ;
			LAYER M4 ;
			RECT 0.120 172.800 17.255 172.920 ;
			LAYER M4 ;
			RECT 0.120 173.304 17.255 173.424 ;
			LAYER M4 ;
			RECT 0.120 173.808 17.255 173.928 ;
			LAYER M4 ;
			RECT 0.120 174.816 17.255 174.936 ;
			LAYER M4 ;
			RECT 0.120 175.320 17.255 175.440 ;
			LAYER M4 ;
			RECT 0.120 175.824 17.255 175.944 ;
			LAYER M4 ;
			RECT 0.120 176.832 17.255 176.952 ;
			LAYER M4 ;
			RECT 0.120 177.336 17.255 177.456 ;
			LAYER M4 ;
			RECT 0.120 177.840 17.255 177.960 ;
			LAYER M4 ;
			RECT 0.120 178.848 17.255 178.968 ;
			LAYER M4 ;
			RECT 0.120 179.352 17.255 179.472 ;
			LAYER M4 ;
			RECT 0.120 179.856 17.255 179.976 ;
			LAYER M4 ;
			RECT 0.120 180.864 17.255 180.984 ;
			LAYER M4 ;
			RECT 0.120 181.368 17.255 181.488 ;
			LAYER M4 ;
			RECT 0.120 181.872 17.255 181.992 ;
			LAYER M4 ;
			RECT 0.120 182.880 17.255 183.000 ;
			LAYER M4 ;
			RECT 0.120 183.384 17.255 183.504 ;
			LAYER M4 ;
			RECT 0.120 183.888 17.255 184.008 ;
			LAYER M4 ;
			RECT 0.120 184.896 17.255 185.016 ;
			LAYER M4 ;
			RECT 0.120 185.400 17.255 185.520 ;
			LAYER M4 ;
			RECT 0.120 185.904 17.255 186.024 ;
			LAYER M4 ;
			RECT 0.120 186.912 17.255 187.032 ;
			LAYER M4 ;
			RECT 0.120 187.416 17.255 187.536 ;
			LAYER M4 ;
			RECT 0.120 187.920 17.255 188.040 ;
			LAYER M4 ;
			RECT 0.120 188.928 17.255 189.048 ;
			LAYER M4 ;
			RECT 0.120 189.432 17.255 189.552 ;
			LAYER M4 ;
			RECT 0.120 189.936 17.255 190.056 ;
			LAYER M4 ;
			RECT 0.120 190.944 17.255 191.064 ;
			LAYER M4 ;
			RECT 0.120 191.448 17.255 191.568 ;
			LAYER M4 ;
			RECT 0.120 191.952 17.255 192.072 ;
			LAYER M4 ;
			RECT 0.120 192.960 17.255 193.080 ;
			LAYER M4 ;
			RECT 0.120 193.464 17.255 193.584 ;
			LAYER M4 ;
			RECT 0.120 193.968 17.255 194.088 ;
			LAYER M4 ;
			RECT 0.120 194.976 17.255 195.096 ;
			LAYER M4 ;
			RECT 0.120 195.480 17.255 195.600 ;
			LAYER M4 ;
			RECT 0.120 195.984 17.255 196.104 ;
			LAYER M4 ;
			RECT 0.120 196.992 17.255 197.112 ;
			LAYER M4 ;
			RECT 0.120 197.496 17.255 197.616 ;
			LAYER M4 ;
			RECT 0.120 198.000 17.255 198.120 ;
			LAYER M4 ;
			RECT 0.120 199.008 17.255 199.128 ;
			LAYER M4 ;
			RECT 0.120 199.512 17.255 199.632 ;
			LAYER M4 ;
			RECT 0.120 200.016 17.255 200.136 ;
			LAYER M4 ;
			RECT 0.120 201.024 17.255 201.144 ;
			LAYER M4 ;
			RECT 0.120 201.528 17.255 201.648 ;
			LAYER M4 ;
			RECT 0.120 202.032 17.255 202.152 ;
			LAYER M4 ;
			RECT 0.120 203.040 17.255 203.160 ;
			LAYER M4 ;
			RECT 0.120 203.544 17.255 203.664 ;
			LAYER M4 ;
			RECT 0.120 204.048 17.255 204.168 ;
			LAYER M4 ;
			RECT 0.120 205.056 17.255 205.176 ;
			LAYER M4 ;
			RECT 0.120 205.560 17.255 205.680 ;
			LAYER M4 ;
			RECT 0.120 206.064 17.255 206.184 ;
			LAYER M4 ;
			RECT 0.120 207.072 17.255 207.192 ;
			LAYER M4 ;
			RECT 0.120 207.576 17.255 207.696 ;
			LAYER M4 ;
			RECT 0.120 208.080 17.255 208.200 ;
			LAYER M4 ;
			RECT 0.120 209.088 17.255 209.208 ;
			LAYER M4 ;
			RECT 0.120 209.592 17.255 209.712 ;
			LAYER M4 ;
			RECT 0.120 210.096 17.255 210.216 ;
			LAYER M4 ;
			RECT 0.120 211.104 17.255 211.224 ;
			LAYER M4 ;
			RECT 0.120 211.608 17.255 211.728 ;
			LAYER M4 ;
			RECT 0.120 212.112 17.255 212.232 ;
			LAYER M4 ;
			RECT 0.120 213.120 17.255 213.240 ;
			LAYER M4 ;
			RECT 0.120 213.624 17.255 213.744 ;
			LAYER M4 ;
			RECT 0.120 214.128 17.255 214.248 ;
			LAYER M4 ;
			RECT 0.120 215.136 17.255 215.256 ;
			LAYER M4 ;
			RECT 0.120 215.640 17.255 215.760 ;
			LAYER M4 ;
			RECT 0.120 216.144 17.255 216.264 ;
			LAYER M4 ;
			RECT 0.120 217.152 17.255 217.272 ;
			LAYER M4 ;
			RECT 0.120 217.656 17.255 217.776 ;
			LAYER M4 ;
			RECT 0.120 218.160 17.255 218.280 ;
			LAYER M4 ;
			RECT 0.120 219.168 17.255 219.288 ;
			LAYER M4 ;
			RECT 0.120 219.672 17.255 219.792 ;
			LAYER M4 ;
			RECT 0.120 220.176 17.255 220.296 ;
			LAYER M4 ;
			RECT 0.120 221.184 17.255 221.304 ;
			LAYER M4 ;
			RECT 0.120 221.688 17.255 221.808 ;
			LAYER M4 ;
			RECT 0.120 222.192 17.255 222.312 ;
			LAYER M4 ;
			RECT 0.120 223.200 17.255 223.320 ;
			LAYER M4 ;
			RECT 0.120 223.704 17.255 223.824 ;
			LAYER M4 ;
			RECT 0.120 224.208 17.255 224.328 ;
			LAYER M4 ;
			RECT 0.120 225.216 17.255 225.336 ;
			LAYER M4 ;
			RECT 0.120 225.720 17.255 225.840 ;
			LAYER M4 ;
			RECT 0.120 226.224 17.255 226.344 ;
			LAYER M4 ;
			RECT 0.120 227.232 17.255 227.352 ;
			LAYER M4 ;
			RECT 0.120 227.736 17.255 227.856 ;
			LAYER M4 ;
			RECT 0.120 228.240 17.255 228.360 ;
			LAYER M4 ;
			RECT 0.120 229.248 17.255 229.368 ;
			LAYER M4 ;
			RECT 0.120 229.752 17.255 229.872 ;
			LAYER M4 ;
			RECT 0.120 230.256 17.255 230.376 ;
			LAYER M4 ;
			RECT 0.120 231.264 17.255 231.384 ;
			LAYER M4 ;
			RECT 0.120 231.768 17.255 231.888 ;
			LAYER M4 ;
			RECT 0.120 232.272 17.255 232.392 ;
			LAYER M4 ;
			RECT 0.120 233.280 17.255 233.400 ;
			LAYER M4 ;
			RECT 0.120 233.784 17.255 233.904 ;
			LAYER M4 ;
			RECT 0.120 234.288 17.255 234.408 ;
			LAYER M4 ;
			RECT 0.120 235.296 17.255 235.416 ;
			LAYER M4 ;
			RECT 0.120 235.800 17.255 235.920 ;
			LAYER M4 ;
			RECT 0.120 236.304 17.255 236.424 ;
			LAYER M4 ;
			RECT 0.120 237.312 17.255 237.432 ;
			LAYER M4 ;
			RECT 0.120 237.816 17.255 237.936 ;
			LAYER M4 ;
			RECT 0.120 238.320 17.255 238.440 ;
			LAYER M4 ;
			RECT 0.120 239.328 17.255 239.448 ;
			LAYER M4 ;
			RECT 0.120 239.832 17.255 239.952 ;
			LAYER M4 ;
			RECT 0.120 240.336 17.255 240.456 ;
			LAYER M4 ;
			RECT 0.120 241.344 17.255 241.464 ;
			LAYER M4 ;
			RECT 0.120 241.848 17.255 241.968 ;
			LAYER M4 ;
			RECT 0.120 242.352 17.255 242.472 ;
			LAYER M4 ;
			RECT 0.120 243.360 17.255 243.480 ;
			LAYER M4 ;
			RECT 0.120 243.864 17.255 243.984 ;
			LAYER M4 ;
			RECT 0.120 244.368 17.255 244.488 ;
			LAYER M4 ;
			RECT 0.120 245.376 17.255 245.496 ;
			LAYER M4 ;
			RECT 0.120 245.880 17.255 246.000 ;
			LAYER M4 ;
			RECT 0.120 246.384 17.255 246.504 ;
			LAYER M4 ;
			RECT 0.120 247.392 17.255 247.512 ;
			LAYER M4 ;
			RECT 0.120 247.896 17.255 248.016 ;
			LAYER M4 ;
			RECT 0.120 248.400 17.255 248.520 ;
			LAYER M4 ;
			RECT 0.120 249.408 17.255 249.528 ;
			LAYER M4 ;
			RECT 0.120 249.912 17.255 250.032 ;
			LAYER M4 ;
			RECT 0.120 250.416 17.255 250.536 ;
			LAYER M4 ;
			RECT 0.120 251.424 17.255 251.544 ;
			LAYER M4 ;
			RECT 0.120 251.928 17.255 252.048 ;
			LAYER M4 ;
			RECT 0.120 252.432 17.255 252.552 ;
			LAYER M4 ;
			RECT 0.120 253.440 17.255 253.560 ;
			LAYER M4 ;
			RECT 0.120 253.944 17.255 254.064 ;
			LAYER M4 ;
			RECT 0.120 254.448 17.255 254.568 ;
			LAYER M4 ;
			RECT 0.120 255.456 17.255 255.576 ;
			LAYER M4 ;
			RECT 0.120 255.960 17.255 256.080 ;
			LAYER M4 ;
			RECT 0.120 256.464 17.255 256.584 ;
			LAYER M4 ;
			RECT 0.120 257.472 17.255 257.592 ;
			LAYER M4 ;
			RECT 0.120 257.976 17.255 258.096 ;
			LAYER M4 ;
			RECT 0.120 258.480 17.255 258.600 ;
			LAYER M4 ;
			RECT 0.120 259.488 17.255 259.608 ;
			LAYER M4 ;
			RECT 0.120 259.992 17.255 260.112 ;
			LAYER M4 ;
			RECT 0.120 260.496 17.255 260.616 ;
			LAYER M4 ;
			RECT 0.120 261.504 17.255 261.624 ;
			LAYER M4 ;
			RECT 0.120 262.008 17.255 262.128 ;
			LAYER M4 ;
			RECT 0.120 262.512 17.255 262.632 ;
			LAYER M4 ;
			RECT 0.120 263.520 17.255 263.640 ;
			LAYER M4 ;
			RECT 0.120 264.024 17.255 264.144 ;
			LAYER M4 ;
			RECT 0.120 264.528 17.255 264.648 ;
			LAYER M4 ;
			RECT 0.120 265.536 17.255 265.656 ;
			LAYER M4 ;
			RECT 0.120 266.040 17.255 266.160 ;
			LAYER M4 ;
			RECT 0.120 266.544 17.255 266.664 ;
			LAYER M4 ;
			RECT 0.120 267.552 17.255 267.672 ;
			LAYER M4 ;
			RECT 0.120 268.056 17.255 268.176 ;
			LAYER M4 ;
			RECT 0.120 268.560 17.255 268.680 ;
			LAYER M4 ;
			RECT 0.120 269.568 17.255 269.688 ;
			LAYER M4 ;
			RECT 0.120 270.072 17.255 270.192 ;
			LAYER M4 ;
			RECT 0.120 270.576 17.255 270.696 ;
			LAYER M4 ;
			RECT 0.120 271.584 17.255 271.704 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 134.600 17.375 134.680 ;
			LAYER M2 ;
			RECT 17.127 134.600 17.375 134.680 ;
			LAYER M3 ;
			RECT 17.127 134.600 17.375 134.680 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081400 LAYER M1 ;
		ANTENNAMAXAREACAR 2.809400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.120400 LAYER M2 ;
		ANTENNAMAXAREACAR 10.990000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.163600 LAYER M3 ;
		ANTENNAMAXAREACAR 30.908400 LAYER M3 ;
	END WEB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 134.408 17.375 134.488 ;
			LAYER M2 ;
			RECT 17.127 134.408 17.375 134.488 ;
			LAYER M3 ;
			RECT 17.127 134.408 17.375 134.488 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100400 LAYER M1 ;
		ANTENNAMAXAREACAR 9.811400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.230600 LAYER M2 ;
		ANTENNAMAXAREACAR 46.438600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.855800 LAYER M3 ;
		ANTENNAMAXAREACAR 215.957000 LAYER M3 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.127 135.560 17.375 135.640 ;
			LAYER M2 ;
			RECT 17.127 135.560 17.375 135.640 ;
			LAYER M3 ;
			RECT 17.127 135.560 17.375 135.640 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100400 LAYER M1 ;
		ANTENNAMAXAREACAR 9.811400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.230600 LAYER M2 ;
		ANTENNAMAXAREACAR 46.438600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.855800 LAYER M3 ;
		ANTENNAMAXAREACAR 215.957000 LAYER M3 ;
	END WTSEL[1]

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 17.375 272.880 ;
		LAYER M2 ;
		RECT 0.000 0.000 17.375 272.880 ;
		LAYER M3 ;
		RECT 0.000 0.000 17.375 272.880 ;
		LAYER M4 ;
		RECT 0.276 272.329 16.975 272.449 ;
		LAYER M4 ;
		RECT 0.300 0.431 16.975 0.551 ;
		LAYER M4 ;
		RECT 0.783 141.880 15.753 141.957 ;
		LAYER M4 ;
		RECT 1.218 134.837 15.753 134.935 ;
		LAYER M4 ;
		RECT 1.218 135.017 15.753 135.115 ;
		LAYER M4 ;
		RECT 1.218 135.197 15.753 135.295 ;
		LAYER M4 ;
		RECT 1.218 135.749 15.753 135.847 ;
		LAYER M4 ;
		RECT 1.218 135.929 15.753 136.027 ;
		LAYER M4 ;
		RECT 1.218 136.109 15.753 136.207 ;
		LAYER M4 ;
		RECT 1.218 136.695 15.753 136.793 ;
		LAYER M4 ;
		RECT 1.218 136.875 15.753 136.973 ;
		LAYER M4 ;
		RECT 1.218 137.055 15.753 137.153 ;
		LAYER M4 ;
		RECT 1.218 137.607 15.753 137.705 ;
		LAYER M4 ;
		RECT 1.218 137.787 15.753 137.885 ;
		LAYER M4 ;
		RECT 1.218 137.967 15.753 138.065 ;
		LAYER M4 ;
		RECT 1.668 133.885 15.753 133.983 ;
		LAYER M4 ;
		RECT 1.668 134.065 15.753 134.163 ;
		LAYER M4 ;
		RECT 1.668 134.245 15.753 134.343 ;
		LAYER M4 ;
		RECT 8.107 1.330 9.089 1.394 ;
		LAYER M4 ;
		RECT 8.107 2.590 9.089 2.654 ;
		LAYER M4 ;
		RECT 8.107 3.346 9.089 3.410 ;
		LAYER M4 ;
		RECT 8.107 4.606 9.089 4.670 ;
		LAYER M4 ;
		RECT 8.107 5.362 9.089 5.426 ;
		LAYER M4 ;
		RECT 8.107 6.622 9.089 6.686 ;
		LAYER M4 ;
		RECT 8.107 7.378 9.089 7.442 ;
		LAYER M4 ;
		RECT 8.107 8.638 9.089 8.702 ;
		LAYER M4 ;
		RECT 8.107 9.394 9.089 9.458 ;
		LAYER M4 ;
		RECT 8.107 10.654 9.089 10.718 ;
		LAYER M4 ;
		RECT 8.107 11.410 9.089 11.474 ;
		LAYER M4 ;
		RECT 8.107 12.670 9.089 12.734 ;
		LAYER M4 ;
		RECT 8.107 13.426 9.089 13.490 ;
		LAYER M4 ;
		RECT 8.107 14.686 9.089 14.750 ;
		LAYER M4 ;
		RECT 8.107 15.442 9.089 15.506 ;
		LAYER M4 ;
		RECT 8.107 16.702 9.089 16.766 ;
		LAYER M4 ;
		RECT 8.107 17.458 9.089 17.522 ;
		LAYER M4 ;
		RECT 8.107 18.718 9.089 18.782 ;
		LAYER M4 ;
		RECT 8.107 19.474 9.089 19.538 ;
		LAYER M4 ;
		RECT 8.107 20.734 9.089 20.798 ;
		LAYER M4 ;
		RECT 8.107 21.490 9.089 21.554 ;
		LAYER M4 ;
		RECT 8.107 22.750 9.089 22.814 ;
		LAYER M4 ;
		RECT 8.107 23.506 9.089 23.570 ;
		LAYER M4 ;
		RECT 8.107 24.766 9.089 24.830 ;
		LAYER M4 ;
		RECT 8.107 25.522 9.089 25.586 ;
		LAYER M4 ;
		RECT 8.107 26.782 9.089 26.846 ;
		LAYER M4 ;
		RECT 8.107 27.538 9.089 27.602 ;
		LAYER M4 ;
		RECT 8.107 28.798 9.089 28.862 ;
		LAYER M4 ;
		RECT 8.107 29.554 9.089 29.618 ;
		LAYER M4 ;
		RECT 8.107 30.814 9.089 30.878 ;
		LAYER M4 ;
		RECT 8.107 31.570 9.089 31.634 ;
		LAYER M4 ;
		RECT 8.107 32.830 9.089 32.894 ;
		LAYER M4 ;
		RECT 8.107 33.586 9.089 33.650 ;
		LAYER M4 ;
		RECT 8.107 34.846 9.089 34.910 ;
		LAYER M4 ;
		RECT 8.107 35.602 9.089 35.666 ;
		LAYER M4 ;
		RECT 8.107 36.862 9.089 36.926 ;
		LAYER M4 ;
		RECT 8.107 37.618 9.089 37.682 ;
		LAYER M4 ;
		RECT 8.107 38.878 9.089 38.942 ;
		LAYER M4 ;
		RECT 8.107 39.634 9.089 39.698 ;
		LAYER M4 ;
		RECT 8.107 40.894 9.089 40.958 ;
		LAYER M4 ;
		RECT 8.107 41.650 9.089 41.714 ;
		LAYER M4 ;
		RECT 8.107 42.910 9.089 42.974 ;
		LAYER M4 ;
		RECT 8.107 43.666 9.089 43.730 ;
		LAYER M4 ;
		RECT 8.107 44.926 9.089 44.990 ;
		LAYER M4 ;
		RECT 8.107 45.682 9.089 45.746 ;
		LAYER M4 ;
		RECT 8.107 46.942 9.089 47.006 ;
		LAYER M4 ;
		RECT 8.107 47.698 9.089 47.762 ;
		LAYER M4 ;
		RECT 8.107 48.958 9.089 49.022 ;
		LAYER M4 ;
		RECT 8.107 49.714 9.089 49.778 ;
		LAYER M4 ;
		RECT 8.107 50.974 9.089 51.038 ;
		LAYER M4 ;
		RECT 8.107 51.730 9.089 51.794 ;
		LAYER M4 ;
		RECT 8.107 52.990 9.089 53.054 ;
		LAYER M4 ;
		RECT 8.107 53.746 9.089 53.810 ;
		LAYER M4 ;
		RECT 8.107 55.006 9.089 55.070 ;
		LAYER M4 ;
		RECT 8.107 55.762 9.089 55.826 ;
		LAYER M4 ;
		RECT 8.107 57.022 9.089 57.086 ;
		LAYER M4 ;
		RECT 8.107 57.778 9.089 57.842 ;
		LAYER M4 ;
		RECT 8.107 59.038 9.089 59.102 ;
		LAYER M4 ;
		RECT 8.107 59.794 9.089 59.858 ;
		LAYER M4 ;
		RECT 8.107 61.054 9.089 61.118 ;
		LAYER M4 ;
		RECT 8.107 61.810 9.089 61.874 ;
		LAYER M4 ;
		RECT 8.107 63.070 9.089 63.134 ;
		LAYER M4 ;
		RECT 8.107 63.826 9.089 63.890 ;
		LAYER M4 ;
		RECT 8.107 65.086 9.089 65.150 ;
		LAYER M4 ;
		RECT 8.107 65.842 9.089 65.906 ;
		LAYER M4 ;
		RECT 8.107 67.102 9.089 67.166 ;
		LAYER M4 ;
		RECT 8.107 67.858 9.089 67.922 ;
		LAYER M4 ;
		RECT 8.107 69.118 9.089 69.182 ;
		LAYER M4 ;
		RECT 8.107 69.874 9.089 69.938 ;
		LAYER M4 ;
		RECT 8.107 71.134 9.089 71.198 ;
		LAYER M4 ;
		RECT 8.107 71.890 9.089 71.954 ;
		LAYER M4 ;
		RECT 8.107 73.150 9.089 73.214 ;
		LAYER M4 ;
		RECT 8.107 73.906 9.089 73.970 ;
		LAYER M4 ;
		RECT 8.107 75.166 9.089 75.230 ;
		LAYER M4 ;
		RECT 8.107 75.922 9.089 75.986 ;
		LAYER M4 ;
		RECT 8.107 77.182 9.089 77.246 ;
		LAYER M4 ;
		RECT 8.107 77.938 9.089 78.002 ;
		LAYER M4 ;
		RECT 8.107 79.198 9.089 79.262 ;
		LAYER M4 ;
		RECT 8.107 79.954 9.089 80.018 ;
		LAYER M4 ;
		RECT 8.107 81.214 9.089 81.278 ;
		LAYER M4 ;
		RECT 8.107 81.970 9.089 82.034 ;
		LAYER M4 ;
		RECT 8.107 83.230 9.089 83.294 ;
		LAYER M4 ;
		RECT 8.107 83.986 9.089 84.050 ;
		LAYER M4 ;
		RECT 8.107 85.246 9.089 85.310 ;
		LAYER M4 ;
		RECT 8.107 86.002 9.089 86.066 ;
		LAYER M4 ;
		RECT 8.107 87.262 9.089 87.326 ;
		LAYER M4 ;
		RECT 8.107 88.018 9.089 88.082 ;
		LAYER M4 ;
		RECT 8.107 89.278 9.089 89.342 ;
		LAYER M4 ;
		RECT 8.107 90.034 9.089 90.098 ;
		LAYER M4 ;
		RECT 8.107 91.294 9.089 91.358 ;
		LAYER M4 ;
		RECT 8.107 92.050 9.089 92.114 ;
		LAYER M4 ;
		RECT 8.107 93.310 9.089 93.374 ;
		LAYER M4 ;
		RECT 8.107 94.066 9.089 94.130 ;
		LAYER M4 ;
		RECT 8.107 95.326 9.089 95.390 ;
		LAYER M4 ;
		RECT 8.107 96.082 9.089 96.146 ;
		LAYER M4 ;
		RECT 8.107 97.342 9.089 97.406 ;
		LAYER M4 ;
		RECT 8.107 98.098 9.089 98.162 ;
		LAYER M4 ;
		RECT 8.107 99.358 9.089 99.422 ;
		LAYER M4 ;
		RECT 8.107 100.114 9.089 100.178 ;
		LAYER M4 ;
		RECT 8.107 101.374 9.089 101.438 ;
		LAYER M4 ;
		RECT 8.107 102.130 9.089 102.194 ;
		LAYER M4 ;
		RECT 8.107 103.390 9.089 103.454 ;
		LAYER M4 ;
		RECT 8.107 104.146 9.089 104.210 ;
		LAYER M4 ;
		RECT 8.107 105.406 9.089 105.470 ;
		LAYER M4 ;
		RECT 8.107 106.162 9.089 106.226 ;
		LAYER M4 ;
		RECT 8.107 107.422 9.089 107.486 ;
		LAYER M4 ;
		RECT 8.107 108.178 9.089 108.242 ;
		LAYER M4 ;
		RECT 8.107 109.438 9.089 109.502 ;
		LAYER M4 ;
		RECT 8.107 110.194 9.089 110.258 ;
		LAYER M4 ;
		RECT 8.107 111.454 9.089 111.518 ;
		LAYER M4 ;
		RECT 8.107 112.210 9.089 112.274 ;
		LAYER M4 ;
		RECT 8.107 113.470 9.089 113.534 ;
		LAYER M4 ;
		RECT 8.107 114.226 9.089 114.290 ;
		LAYER M4 ;
		RECT 8.107 115.486 9.089 115.550 ;
		LAYER M4 ;
		RECT 8.107 116.242 9.089 116.306 ;
		LAYER M4 ;
		RECT 8.107 117.502 9.089 117.566 ;
		LAYER M4 ;
		RECT 8.107 118.258 9.089 118.322 ;
		LAYER M4 ;
		RECT 8.107 119.518 9.089 119.582 ;
		LAYER M4 ;
		RECT 8.107 120.274 9.089 120.338 ;
		LAYER M4 ;
		RECT 8.107 121.534 9.089 121.598 ;
		LAYER M4 ;
		RECT 8.107 122.290 9.089 122.354 ;
		LAYER M4 ;
		RECT 8.107 123.550 9.089 123.614 ;
		LAYER M4 ;
		RECT 8.107 124.306 9.089 124.370 ;
		LAYER M4 ;
		RECT 8.107 125.566 9.089 125.630 ;
		LAYER M4 ;
		RECT 8.107 126.322 9.089 126.386 ;
		LAYER M4 ;
		RECT 8.107 127.582 9.089 127.646 ;
		LAYER M4 ;
		RECT 8.107 128.338 9.089 128.402 ;
		LAYER M4 ;
		RECT 8.107 129.598 9.089 129.662 ;
		LAYER M4 ;
		RECT 8.107 143.218 9.089 143.282 ;
		LAYER M4 ;
		RECT 8.107 144.478 9.089 144.542 ;
		LAYER M4 ;
		RECT 8.107 145.234 9.089 145.298 ;
		LAYER M4 ;
		RECT 8.107 146.494 9.089 146.558 ;
		LAYER M4 ;
		RECT 8.107 147.250 9.089 147.314 ;
		LAYER M4 ;
		RECT 8.107 148.510 9.089 148.574 ;
		LAYER M4 ;
		RECT 8.107 149.266 9.089 149.330 ;
		LAYER M4 ;
		RECT 8.107 150.526 9.089 150.590 ;
		LAYER M4 ;
		RECT 8.107 151.282 9.089 151.346 ;
		LAYER M4 ;
		RECT 8.107 152.542 9.089 152.606 ;
		LAYER M4 ;
		RECT 8.107 153.298 9.089 153.362 ;
		LAYER M4 ;
		RECT 8.107 154.558 9.089 154.622 ;
		LAYER M4 ;
		RECT 8.107 155.314 9.089 155.378 ;
		LAYER M4 ;
		RECT 8.107 156.574 9.089 156.638 ;
		LAYER M4 ;
		RECT 8.107 157.330 9.089 157.394 ;
		LAYER M4 ;
		RECT 8.107 158.590 9.089 158.654 ;
		LAYER M4 ;
		RECT 8.107 159.346 9.089 159.410 ;
		LAYER M4 ;
		RECT 8.107 160.606 9.089 160.670 ;
		LAYER M4 ;
		RECT 8.107 161.362 9.089 161.426 ;
		LAYER M4 ;
		RECT 8.107 162.622 9.089 162.686 ;
		LAYER M4 ;
		RECT 8.107 163.378 9.089 163.442 ;
		LAYER M4 ;
		RECT 8.107 164.638 9.089 164.702 ;
		LAYER M4 ;
		RECT 8.107 165.394 9.089 165.458 ;
		LAYER M4 ;
		RECT 8.107 166.654 9.089 166.718 ;
		LAYER M4 ;
		RECT 8.107 167.410 9.089 167.474 ;
		LAYER M4 ;
		RECT 8.107 168.670 9.089 168.734 ;
		LAYER M4 ;
		RECT 8.107 169.426 9.089 169.490 ;
		LAYER M4 ;
		RECT 8.107 170.686 9.089 170.750 ;
		LAYER M4 ;
		RECT 8.107 171.442 9.089 171.506 ;
		LAYER M4 ;
		RECT 8.107 172.702 9.089 172.766 ;
		LAYER M4 ;
		RECT 8.107 173.458 9.089 173.522 ;
		LAYER M4 ;
		RECT 8.107 174.718 9.089 174.782 ;
		LAYER M4 ;
		RECT 8.107 175.474 9.089 175.538 ;
		LAYER M4 ;
		RECT 8.107 176.734 9.089 176.798 ;
		LAYER M4 ;
		RECT 8.107 177.490 9.089 177.554 ;
		LAYER M4 ;
		RECT 8.107 178.750 9.089 178.814 ;
		LAYER M4 ;
		RECT 8.107 179.506 9.089 179.570 ;
		LAYER M4 ;
		RECT 8.107 180.766 9.089 180.830 ;
		LAYER M4 ;
		RECT 8.107 181.522 9.089 181.586 ;
		LAYER M4 ;
		RECT 8.107 182.782 9.089 182.846 ;
		LAYER M4 ;
		RECT 8.107 183.538 9.089 183.602 ;
		LAYER M4 ;
		RECT 8.107 184.798 9.089 184.862 ;
		LAYER M4 ;
		RECT 8.107 185.554 9.089 185.618 ;
		LAYER M4 ;
		RECT 8.107 186.814 9.089 186.878 ;
		LAYER M4 ;
		RECT 8.107 187.570 9.089 187.634 ;
		LAYER M4 ;
		RECT 8.107 188.830 9.089 188.894 ;
		LAYER M4 ;
		RECT 8.107 189.586 9.089 189.650 ;
		LAYER M4 ;
		RECT 8.107 190.846 9.089 190.910 ;
		LAYER M4 ;
		RECT 8.107 191.602 9.089 191.666 ;
		LAYER M4 ;
		RECT 8.107 192.862 9.089 192.926 ;
		LAYER M4 ;
		RECT 8.107 193.618 9.089 193.682 ;
		LAYER M4 ;
		RECT 8.107 194.878 9.089 194.942 ;
		LAYER M4 ;
		RECT 8.107 195.634 9.089 195.698 ;
		LAYER M4 ;
		RECT 8.107 196.894 9.089 196.958 ;
		LAYER M4 ;
		RECT 8.107 197.650 9.089 197.714 ;
		LAYER M4 ;
		RECT 8.107 198.910 9.089 198.974 ;
		LAYER M4 ;
		RECT 8.107 199.666 9.089 199.730 ;
		LAYER M4 ;
		RECT 8.107 200.926 9.089 200.990 ;
		LAYER M4 ;
		RECT 8.107 201.682 9.089 201.746 ;
		LAYER M4 ;
		RECT 8.107 202.942 9.089 203.006 ;
		LAYER M4 ;
		RECT 8.107 203.698 9.089 203.762 ;
		LAYER M4 ;
		RECT 8.107 204.958 9.089 205.022 ;
		LAYER M4 ;
		RECT 8.107 205.714 9.089 205.778 ;
		LAYER M4 ;
		RECT 8.107 206.974 9.089 207.038 ;
		LAYER M4 ;
		RECT 8.107 207.730 9.089 207.794 ;
		LAYER M4 ;
		RECT 8.107 208.990 9.089 209.054 ;
		LAYER M4 ;
		RECT 8.107 209.746 9.089 209.810 ;
		LAYER M4 ;
		RECT 8.107 211.006 9.089 211.070 ;
		LAYER M4 ;
		RECT 8.107 211.762 9.089 211.826 ;
		LAYER M4 ;
		RECT 8.107 213.022 9.089 213.086 ;
		LAYER M4 ;
		RECT 8.107 213.778 9.089 213.842 ;
		LAYER M4 ;
		RECT 8.107 215.038 9.089 215.102 ;
		LAYER M4 ;
		RECT 8.107 215.794 9.089 215.858 ;
		LAYER M4 ;
		RECT 8.107 217.054 9.089 217.118 ;
		LAYER M4 ;
		RECT 8.107 217.810 9.089 217.874 ;
		LAYER M4 ;
		RECT 8.107 219.070 9.089 219.134 ;
		LAYER M4 ;
		RECT 8.107 219.826 9.089 219.890 ;
		LAYER M4 ;
		RECT 8.107 221.086 9.089 221.150 ;
		LAYER M4 ;
		RECT 8.107 221.842 9.089 221.906 ;
		LAYER M4 ;
		RECT 8.107 223.102 9.089 223.166 ;
		LAYER M4 ;
		RECT 8.107 223.858 9.089 223.922 ;
		LAYER M4 ;
		RECT 8.107 225.118 9.089 225.182 ;
		LAYER M4 ;
		RECT 8.107 225.874 9.089 225.938 ;
		LAYER M4 ;
		RECT 8.107 227.134 9.089 227.198 ;
		LAYER M4 ;
		RECT 8.107 227.890 9.089 227.954 ;
		LAYER M4 ;
		RECT 8.107 229.150 9.089 229.214 ;
		LAYER M4 ;
		RECT 8.107 229.906 9.089 229.970 ;
		LAYER M4 ;
		RECT 8.107 231.166 9.089 231.230 ;
		LAYER M4 ;
		RECT 8.107 231.922 9.089 231.986 ;
		LAYER M4 ;
		RECT 8.107 233.182 9.089 233.246 ;
		LAYER M4 ;
		RECT 8.107 233.938 9.089 234.002 ;
		LAYER M4 ;
		RECT 8.107 235.198 9.089 235.262 ;
		LAYER M4 ;
		RECT 8.107 235.954 9.089 236.018 ;
		LAYER M4 ;
		RECT 8.107 237.214 9.089 237.278 ;
		LAYER M4 ;
		RECT 8.107 237.970 9.089 238.034 ;
		LAYER M4 ;
		RECT 8.107 239.230 9.089 239.294 ;
		LAYER M4 ;
		RECT 8.107 239.986 9.089 240.050 ;
		LAYER M4 ;
		RECT 8.107 241.246 9.089 241.310 ;
		LAYER M4 ;
		RECT 8.107 242.002 9.089 242.066 ;
		LAYER M4 ;
		RECT 8.107 243.262 9.089 243.326 ;
		LAYER M4 ;
		RECT 8.107 244.018 9.089 244.082 ;
		LAYER M4 ;
		RECT 8.107 245.278 9.089 245.342 ;
		LAYER M4 ;
		RECT 8.107 246.034 9.089 246.098 ;
		LAYER M4 ;
		RECT 8.107 247.294 9.089 247.358 ;
		LAYER M4 ;
		RECT 8.107 248.050 9.089 248.114 ;
		LAYER M4 ;
		RECT 8.107 249.310 9.089 249.374 ;
		LAYER M4 ;
		RECT 8.107 250.066 9.089 250.130 ;
		LAYER M4 ;
		RECT 8.107 251.326 9.089 251.390 ;
		LAYER M4 ;
		RECT 8.107 252.082 9.089 252.146 ;
		LAYER M4 ;
		RECT 8.107 253.342 9.089 253.406 ;
		LAYER M4 ;
		RECT 8.107 254.098 9.089 254.162 ;
		LAYER M4 ;
		RECT 8.107 255.358 9.089 255.422 ;
		LAYER M4 ;
		RECT 8.107 256.114 9.089 256.178 ;
		LAYER M4 ;
		RECT 8.107 257.374 9.089 257.438 ;
		LAYER M4 ;
		RECT 8.107 258.130 9.089 258.194 ;
		LAYER M4 ;
		RECT 8.107 259.390 9.089 259.454 ;
		LAYER M4 ;
		RECT 8.107 260.146 9.089 260.210 ;
		LAYER M4 ;
		RECT 8.107 261.406 9.089 261.470 ;
		LAYER M4 ;
		RECT 8.107 262.162 9.089 262.226 ;
		LAYER M4 ;
		RECT 8.107 263.422 9.089 263.486 ;
		LAYER M4 ;
		RECT 8.107 264.178 9.089 264.242 ;
		LAYER M4 ;
		RECT 8.107 265.438 9.089 265.502 ;
		LAYER M4 ;
		RECT 8.107 266.194 9.089 266.258 ;
		LAYER M4 ;
		RECT 8.107 267.454 9.089 267.518 ;
		LAYER M4 ;
		RECT 8.107 268.210 9.089 268.274 ;
		LAYER M4 ;
		RECT 8.107 269.470 9.089 269.534 ;
		LAYER M4 ;
		RECT 8.107 270.226 9.089 270.290 ;
		LAYER M4 ;
		RECT 8.107 271.486 9.089 271.550 ;
		LAYER M4 ;
		RECT 9.616 1.337 11.339 1.387 ;
		LAYER M4 ;
		RECT 9.616 2.597 11.531 2.647 ;
		LAYER M4 ;
		RECT 9.616 3.353 11.339 3.403 ;
		LAYER M4 ;
		RECT 9.616 4.613 11.531 4.663 ;
		LAYER M4 ;
		RECT 9.616 5.369 11.339 5.419 ;
		LAYER M4 ;
		RECT 9.616 6.629 11.531 6.679 ;
		LAYER M4 ;
		RECT 9.616 7.385 11.339 7.435 ;
		LAYER M4 ;
		RECT 9.616 8.645 11.531 8.695 ;
		LAYER M4 ;
		RECT 9.616 9.401 11.339 9.451 ;
		LAYER M4 ;
		RECT 9.616 10.661 11.531 10.711 ;
		LAYER M4 ;
		RECT 9.616 11.417 11.339 11.467 ;
		LAYER M4 ;
		RECT 9.616 12.677 11.531 12.727 ;
		LAYER M4 ;
		RECT 9.616 13.433 11.339 13.483 ;
		LAYER M4 ;
		RECT 9.616 14.693 11.531 14.743 ;
		LAYER M4 ;
		RECT 9.616 15.449 11.339 15.499 ;
		LAYER M4 ;
		RECT 9.616 16.709 11.531 16.759 ;
		LAYER M4 ;
		RECT 9.616 17.465 11.339 17.515 ;
		LAYER M4 ;
		RECT 9.616 18.725 11.531 18.775 ;
		LAYER M4 ;
		RECT 9.616 19.481 11.339 19.531 ;
		LAYER M4 ;
		RECT 9.616 20.741 11.531 20.791 ;
		LAYER M4 ;
		RECT 9.616 21.497 11.339 21.547 ;
		LAYER M4 ;
		RECT 9.616 22.757 11.531 22.807 ;
		LAYER M4 ;
		RECT 9.616 23.513 11.339 23.563 ;
		LAYER M4 ;
		RECT 9.616 24.773 11.531 24.823 ;
		LAYER M4 ;
		RECT 9.616 25.529 11.339 25.579 ;
		LAYER M4 ;
		RECT 9.616 26.789 11.531 26.839 ;
		LAYER M4 ;
		RECT 9.616 27.545 11.339 27.595 ;
		LAYER M4 ;
		RECT 9.616 28.805 11.531 28.855 ;
		LAYER M4 ;
		RECT 9.616 29.561 11.339 29.611 ;
		LAYER M4 ;
		RECT 9.616 30.821 11.531 30.871 ;
		LAYER M4 ;
		RECT 9.616 31.577 11.339 31.627 ;
		LAYER M4 ;
		RECT 9.616 32.837 11.531 32.887 ;
		LAYER M4 ;
		RECT 9.616 33.593 11.339 33.643 ;
		LAYER M4 ;
		RECT 9.616 34.853 11.531 34.903 ;
		LAYER M4 ;
		RECT 9.616 35.609 11.339 35.659 ;
		LAYER M4 ;
		RECT 9.616 36.869 11.531 36.919 ;
		LAYER M4 ;
		RECT 9.616 37.625 11.339 37.675 ;
		LAYER M4 ;
		RECT 9.616 38.885 11.531 38.935 ;
		LAYER M4 ;
		RECT 9.616 39.641 11.339 39.691 ;
		LAYER M4 ;
		RECT 9.616 40.901 11.531 40.951 ;
		LAYER M4 ;
		RECT 9.616 41.657 11.339 41.707 ;
		LAYER M4 ;
		RECT 9.616 42.917 11.531 42.967 ;
		LAYER M4 ;
		RECT 9.616 43.673 11.339 43.723 ;
		LAYER M4 ;
		RECT 9.616 44.933 11.531 44.983 ;
		LAYER M4 ;
		RECT 9.616 45.689 11.339 45.739 ;
		LAYER M4 ;
		RECT 9.616 46.949 11.531 46.999 ;
		LAYER M4 ;
		RECT 9.616 47.705 11.339 47.755 ;
		LAYER M4 ;
		RECT 9.616 48.965 11.531 49.015 ;
		LAYER M4 ;
		RECT 9.616 49.721 11.339 49.771 ;
		LAYER M4 ;
		RECT 9.616 50.981 11.531 51.031 ;
		LAYER M4 ;
		RECT 9.616 51.737 11.339 51.787 ;
		LAYER M4 ;
		RECT 9.616 52.997 11.531 53.047 ;
		LAYER M4 ;
		RECT 9.616 53.753 11.339 53.803 ;
		LAYER M4 ;
		RECT 9.616 55.013 11.531 55.063 ;
		LAYER M4 ;
		RECT 9.616 55.769 11.339 55.819 ;
		LAYER M4 ;
		RECT 9.616 57.029 11.531 57.079 ;
		LAYER M4 ;
		RECT 9.616 57.785 11.339 57.835 ;
		LAYER M4 ;
		RECT 9.616 59.045 11.531 59.095 ;
		LAYER M4 ;
		RECT 9.616 59.801 11.339 59.851 ;
		LAYER M4 ;
		RECT 9.616 61.061 11.531 61.111 ;
		LAYER M4 ;
		RECT 9.616 61.817 11.339 61.867 ;
		LAYER M4 ;
		RECT 9.616 63.077 11.531 63.127 ;
		LAYER M4 ;
		RECT 9.616 63.833 11.339 63.883 ;
		LAYER M4 ;
		RECT 9.616 65.093 11.531 65.143 ;
		LAYER M4 ;
		RECT 9.616 65.849 11.339 65.899 ;
		LAYER M4 ;
		RECT 9.616 67.109 11.531 67.159 ;
		LAYER M4 ;
		RECT 9.616 67.865 11.339 67.915 ;
		LAYER M4 ;
		RECT 9.616 69.125 11.531 69.175 ;
		LAYER M4 ;
		RECT 9.616 69.881 11.339 69.931 ;
		LAYER M4 ;
		RECT 9.616 71.141 11.531 71.191 ;
		LAYER M4 ;
		RECT 9.616 71.897 11.339 71.947 ;
		LAYER M4 ;
		RECT 9.616 73.157 11.531 73.207 ;
		LAYER M4 ;
		RECT 9.616 73.913 11.339 73.963 ;
		LAYER M4 ;
		RECT 9.616 75.173 11.531 75.223 ;
		LAYER M4 ;
		RECT 9.616 75.929 11.339 75.979 ;
		LAYER M4 ;
		RECT 9.616 77.189 11.531 77.239 ;
		LAYER M4 ;
		RECT 9.616 77.945 11.339 77.995 ;
		LAYER M4 ;
		RECT 9.616 79.205 11.531 79.255 ;
		LAYER M4 ;
		RECT 9.616 79.961 11.339 80.011 ;
		LAYER M4 ;
		RECT 9.616 81.221 11.531 81.271 ;
		LAYER M4 ;
		RECT 9.616 81.977 11.339 82.027 ;
		LAYER M4 ;
		RECT 9.616 83.237 11.531 83.287 ;
		LAYER M4 ;
		RECT 9.616 83.993 11.339 84.043 ;
		LAYER M4 ;
		RECT 9.616 85.253 11.531 85.303 ;
		LAYER M4 ;
		RECT 9.616 86.009 11.339 86.059 ;
		LAYER M4 ;
		RECT 9.616 87.269 11.531 87.319 ;
		LAYER M4 ;
		RECT 9.616 88.025 11.339 88.075 ;
		LAYER M4 ;
		RECT 9.616 89.285 11.531 89.335 ;
		LAYER M4 ;
		RECT 9.616 90.041 11.339 90.091 ;
		LAYER M4 ;
		RECT 9.616 91.301 11.531 91.351 ;
		LAYER M4 ;
		RECT 9.616 92.057 11.339 92.107 ;
		LAYER M4 ;
		RECT 9.616 93.317 11.531 93.367 ;
		LAYER M4 ;
		RECT 9.616 94.073 11.339 94.123 ;
		LAYER M4 ;
		RECT 9.616 95.333 11.531 95.383 ;
		LAYER M4 ;
		RECT 9.616 96.089 11.339 96.139 ;
		LAYER M4 ;
		RECT 9.616 97.349 11.531 97.399 ;
		LAYER M4 ;
		RECT 9.616 98.105 11.339 98.155 ;
		LAYER M4 ;
		RECT 9.616 99.365 11.531 99.415 ;
		LAYER M4 ;
		RECT 9.616 100.121 11.339 100.171 ;
		LAYER M4 ;
		RECT 9.616 101.381 11.531 101.431 ;
		LAYER M4 ;
		RECT 9.616 102.137 11.339 102.187 ;
		LAYER M4 ;
		RECT 9.616 103.397 11.531 103.447 ;
		LAYER M4 ;
		RECT 9.616 104.153 11.339 104.203 ;
		LAYER M4 ;
		RECT 9.616 105.413 11.531 105.463 ;
		LAYER M4 ;
		RECT 9.616 106.169 11.339 106.219 ;
		LAYER M4 ;
		RECT 9.616 107.429 11.531 107.479 ;
		LAYER M4 ;
		RECT 9.616 108.185 11.339 108.235 ;
		LAYER M4 ;
		RECT 9.616 109.445 11.531 109.495 ;
		LAYER M4 ;
		RECT 9.616 110.201 11.339 110.251 ;
		LAYER M4 ;
		RECT 9.616 111.461 11.531 111.511 ;
		LAYER M4 ;
		RECT 9.616 112.217 11.339 112.267 ;
		LAYER M4 ;
		RECT 9.616 113.477 11.531 113.527 ;
		LAYER M4 ;
		RECT 9.616 114.233 11.339 114.283 ;
		LAYER M4 ;
		RECT 9.616 115.493 11.531 115.543 ;
		LAYER M4 ;
		RECT 9.616 116.249 11.339 116.299 ;
		LAYER M4 ;
		RECT 9.616 117.509 11.531 117.559 ;
		LAYER M4 ;
		RECT 9.616 118.265 11.339 118.315 ;
		LAYER M4 ;
		RECT 9.616 119.525 11.531 119.575 ;
		LAYER M4 ;
		RECT 9.616 120.281 11.339 120.331 ;
		LAYER M4 ;
		RECT 9.616 121.541 11.531 121.591 ;
		LAYER M4 ;
		RECT 9.616 122.297 11.339 122.347 ;
		LAYER M4 ;
		RECT 9.616 123.557 11.531 123.607 ;
		LAYER M4 ;
		RECT 9.616 124.313 11.339 124.363 ;
		LAYER M4 ;
		RECT 9.616 125.573 11.531 125.623 ;
		LAYER M4 ;
		RECT 9.616 126.329 11.339 126.379 ;
		LAYER M4 ;
		RECT 9.616 127.589 11.531 127.639 ;
		LAYER M4 ;
		RECT 9.616 128.345 11.339 128.395 ;
		LAYER M4 ;
		RECT 9.616 129.605 11.531 129.655 ;
		LAYER M4 ;
		RECT 9.616 143.225 11.339 143.275 ;
		LAYER M4 ;
		RECT 9.616 144.485 11.531 144.535 ;
		LAYER M4 ;
		RECT 9.616 145.241 11.339 145.291 ;
		LAYER M4 ;
		RECT 9.616 146.501 11.531 146.551 ;
		LAYER M4 ;
		RECT 9.616 147.257 11.339 147.307 ;
		LAYER M4 ;
		RECT 9.616 148.517 11.531 148.567 ;
		LAYER M4 ;
		RECT 9.616 149.273 11.339 149.323 ;
		LAYER M4 ;
		RECT 9.616 150.533 11.531 150.583 ;
		LAYER M4 ;
		RECT 9.616 151.289 11.339 151.339 ;
		LAYER M4 ;
		RECT 9.616 152.549 11.531 152.599 ;
		LAYER M4 ;
		RECT 9.616 153.305 11.339 153.355 ;
		LAYER M4 ;
		RECT 9.616 154.565 11.531 154.615 ;
		LAYER M4 ;
		RECT 9.616 155.321 11.339 155.371 ;
		LAYER M4 ;
		RECT 9.616 156.581 11.531 156.631 ;
		LAYER M4 ;
		RECT 9.616 157.337 11.339 157.387 ;
		LAYER M4 ;
		RECT 9.616 158.597 11.531 158.647 ;
		LAYER M4 ;
		RECT 9.616 159.353 11.339 159.403 ;
		LAYER M4 ;
		RECT 9.616 160.613 11.531 160.663 ;
		LAYER M4 ;
		RECT 9.616 161.369 11.339 161.419 ;
		LAYER M4 ;
		RECT 9.616 162.629 11.531 162.679 ;
		LAYER M4 ;
		RECT 9.616 163.385 11.339 163.435 ;
		LAYER M4 ;
		RECT 9.616 164.645 11.531 164.695 ;
		LAYER M4 ;
		RECT 9.616 165.401 11.339 165.451 ;
		LAYER M4 ;
		RECT 9.616 166.661 11.531 166.711 ;
		LAYER M4 ;
		RECT 9.616 167.417 11.339 167.467 ;
		LAYER M4 ;
		RECT 9.616 168.677 11.531 168.727 ;
		LAYER M4 ;
		RECT 9.616 169.433 11.339 169.483 ;
		LAYER M4 ;
		RECT 9.616 170.693 11.531 170.743 ;
		LAYER M4 ;
		RECT 9.616 171.449 11.339 171.499 ;
		LAYER M4 ;
		RECT 9.616 172.709 11.531 172.759 ;
		LAYER M4 ;
		RECT 9.616 173.465 11.339 173.515 ;
		LAYER M4 ;
		RECT 9.616 174.725 11.531 174.775 ;
		LAYER M4 ;
		RECT 9.616 175.481 11.339 175.531 ;
		LAYER M4 ;
		RECT 9.616 176.741 11.531 176.791 ;
		LAYER M4 ;
		RECT 9.616 177.497 11.339 177.547 ;
		LAYER M4 ;
		RECT 9.616 178.757 11.531 178.807 ;
		LAYER M4 ;
		RECT 9.616 179.513 11.339 179.563 ;
		LAYER M4 ;
		RECT 9.616 180.773 11.531 180.823 ;
		LAYER M4 ;
		RECT 9.616 181.529 11.339 181.579 ;
		LAYER M4 ;
		RECT 9.616 182.789 11.531 182.839 ;
		LAYER M4 ;
		RECT 9.616 183.545 11.339 183.595 ;
		LAYER M4 ;
		RECT 9.616 184.805 11.531 184.855 ;
		LAYER M4 ;
		RECT 9.616 185.561 11.339 185.611 ;
		LAYER M4 ;
		RECT 9.616 186.821 11.531 186.871 ;
		LAYER M4 ;
		RECT 9.616 187.577 11.339 187.627 ;
		LAYER M4 ;
		RECT 9.616 188.837 11.531 188.887 ;
		LAYER M4 ;
		RECT 9.616 189.593 11.339 189.643 ;
		LAYER M4 ;
		RECT 9.616 190.853 11.531 190.903 ;
		LAYER M4 ;
		RECT 9.616 191.609 11.339 191.659 ;
		LAYER M4 ;
		RECT 9.616 192.869 11.531 192.919 ;
		LAYER M4 ;
		RECT 9.616 193.625 11.339 193.675 ;
		LAYER M4 ;
		RECT 9.616 194.885 11.531 194.935 ;
		LAYER M4 ;
		RECT 9.616 195.641 11.339 195.691 ;
		LAYER M4 ;
		RECT 9.616 196.901 11.531 196.951 ;
		LAYER M4 ;
		RECT 9.616 197.657 11.339 197.707 ;
		LAYER M4 ;
		RECT 9.616 198.917 11.531 198.967 ;
		LAYER M4 ;
		RECT 9.616 199.673 11.339 199.723 ;
		LAYER M4 ;
		RECT 9.616 200.933 11.531 200.983 ;
		LAYER M4 ;
		RECT 9.616 201.689 11.339 201.739 ;
		LAYER M4 ;
		RECT 9.616 202.949 11.531 202.999 ;
		LAYER M4 ;
		RECT 9.616 203.705 11.339 203.755 ;
		LAYER M4 ;
		RECT 9.616 204.965 11.531 205.015 ;
		LAYER M4 ;
		RECT 9.616 205.721 11.339 205.771 ;
		LAYER M4 ;
		RECT 9.616 206.981 11.531 207.031 ;
		LAYER M4 ;
		RECT 9.616 207.737 11.339 207.787 ;
		LAYER M4 ;
		RECT 9.616 208.997 11.531 209.047 ;
		LAYER M4 ;
		RECT 9.616 209.753 11.339 209.803 ;
		LAYER M4 ;
		RECT 9.616 211.013 11.531 211.063 ;
		LAYER M4 ;
		RECT 9.616 211.769 11.339 211.819 ;
		LAYER M4 ;
		RECT 9.616 213.029 11.531 213.079 ;
		LAYER M4 ;
		RECT 9.616 213.785 11.339 213.835 ;
		LAYER M4 ;
		RECT 9.616 215.045 11.531 215.095 ;
		LAYER M4 ;
		RECT 9.616 215.801 11.339 215.851 ;
		LAYER M4 ;
		RECT 9.616 217.061 11.531 217.111 ;
		LAYER M4 ;
		RECT 9.616 217.817 11.339 217.867 ;
		LAYER M4 ;
		RECT 9.616 219.077 11.531 219.127 ;
		LAYER M4 ;
		RECT 9.616 219.833 11.339 219.883 ;
		LAYER M4 ;
		RECT 9.616 221.093 11.531 221.143 ;
		LAYER M4 ;
		RECT 9.616 221.849 11.339 221.899 ;
		LAYER M4 ;
		RECT 9.616 223.109 11.531 223.159 ;
		LAYER M4 ;
		RECT 9.616 223.865 11.339 223.915 ;
		LAYER M4 ;
		RECT 9.616 225.125 11.531 225.175 ;
		LAYER M4 ;
		RECT 9.616 225.881 11.339 225.931 ;
		LAYER M4 ;
		RECT 9.616 227.141 11.531 227.191 ;
		LAYER M4 ;
		RECT 9.616 227.897 11.339 227.947 ;
		LAYER M4 ;
		RECT 9.616 229.157 11.531 229.207 ;
		LAYER M4 ;
		RECT 9.616 229.913 11.339 229.963 ;
		LAYER M4 ;
		RECT 9.616 231.173 11.531 231.223 ;
		LAYER M4 ;
		RECT 9.616 231.929 11.339 231.979 ;
		LAYER M4 ;
		RECT 9.616 233.189 11.531 233.239 ;
		LAYER M4 ;
		RECT 9.616 233.945 11.339 233.995 ;
		LAYER M4 ;
		RECT 9.616 235.205 11.531 235.255 ;
		LAYER M4 ;
		RECT 9.616 235.961 11.339 236.011 ;
		LAYER M4 ;
		RECT 9.616 237.221 11.531 237.271 ;
		LAYER M4 ;
		RECT 9.616 237.977 11.339 238.027 ;
		LAYER M4 ;
		RECT 9.616 239.237 11.531 239.287 ;
		LAYER M4 ;
		RECT 9.616 239.993 11.339 240.043 ;
		LAYER M4 ;
		RECT 9.616 241.253 11.531 241.303 ;
		LAYER M4 ;
		RECT 9.616 242.009 11.339 242.059 ;
		LAYER M4 ;
		RECT 9.616 243.269 11.531 243.319 ;
		LAYER M4 ;
		RECT 9.616 244.025 11.339 244.075 ;
		LAYER M4 ;
		RECT 9.616 245.285 11.531 245.335 ;
		LAYER M4 ;
		RECT 9.616 246.041 11.339 246.091 ;
		LAYER M4 ;
		RECT 9.616 247.301 11.531 247.351 ;
		LAYER M4 ;
		RECT 9.616 248.057 11.339 248.107 ;
		LAYER M4 ;
		RECT 9.616 249.317 11.531 249.367 ;
		LAYER M4 ;
		RECT 9.616 250.073 11.339 250.123 ;
		LAYER M4 ;
		RECT 9.616 251.333 11.531 251.383 ;
		LAYER M4 ;
		RECT 9.616 252.089 11.339 252.139 ;
		LAYER M4 ;
		RECT 9.616 253.349 11.531 253.399 ;
		LAYER M4 ;
		RECT 9.616 254.105 11.339 254.155 ;
		LAYER M4 ;
		RECT 9.616 255.365 11.531 255.415 ;
		LAYER M4 ;
		RECT 9.616 256.121 11.339 256.171 ;
		LAYER M4 ;
		RECT 9.616 257.381 11.531 257.431 ;
		LAYER M4 ;
		RECT 9.616 258.137 11.339 258.187 ;
		LAYER M4 ;
		RECT 9.616 259.397 11.531 259.447 ;
		LAYER M4 ;
		RECT 9.616 260.153 11.339 260.203 ;
		LAYER M4 ;
		RECT 9.616 261.413 11.531 261.463 ;
		LAYER M4 ;
		RECT 9.616 262.169 11.339 262.219 ;
		LAYER M4 ;
		RECT 9.616 263.429 11.531 263.479 ;
		LAYER M4 ;
		RECT 9.616 264.185 11.339 264.235 ;
		LAYER M4 ;
		RECT 9.616 265.445 11.531 265.495 ;
		LAYER M4 ;
		RECT 9.616 266.201 11.339 266.251 ;
		LAYER M4 ;
		RECT 9.616 267.461 11.531 267.511 ;
		LAYER M4 ;
		RECT 9.616 268.217 11.339 268.267 ;
		LAYER M4 ;
		RECT 9.616 269.477 11.531 269.527 ;
		LAYER M4 ;
		RECT 9.616 270.233 11.339 270.283 ;
		LAYER M4 ;
		RECT 9.616 271.493 11.531 271.543 ;
		LAYER M4 ;
		RECT 10.717 1.589 11.609 1.639 ;
		LAYER M4 ;
		RECT 10.717 2.345 11.609 2.395 ;
		LAYER M4 ;
		RECT 10.717 3.605 11.609 3.655 ;
		LAYER M4 ;
		RECT 10.717 4.361 11.609 4.411 ;
		LAYER M4 ;
		RECT 10.717 5.621 11.609 5.671 ;
		LAYER M4 ;
		RECT 10.717 6.377 11.609 6.427 ;
		LAYER M4 ;
		RECT 10.717 7.637 11.609 7.687 ;
		LAYER M4 ;
		RECT 10.717 8.393 11.609 8.443 ;
		LAYER M4 ;
		RECT 10.717 9.653 11.609 9.703 ;
		LAYER M4 ;
		RECT 10.717 10.409 11.609 10.459 ;
		LAYER M4 ;
		RECT 10.717 11.669 11.609 11.719 ;
		LAYER M4 ;
		RECT 10.717 12.425 11.609 12.475 ;
		LAYER M4 ;
		RECT 10.717 13.685 11.609 13.735 ;
		LAYER M4 ;
		RECT 10.717 14.441 11.609 14.491 ;
		LAYER M4 ;
		RECT 10.717 15.701 11.609 15.751 ;
		LAYER M4 ;
		RECT 10.717 16.457 11.609 16.507 ;
		LAYER M4 ;
		RECT 10.717 17.717 11.609 17.767 ;
		LAYER M4 ;
		RECT 10.717 18.473 11.609 18.523 ;
		LAYER M4 ;
		RECT 10.717 19.733 11.609 19.783 ;
		LAYER M4 ;
		RECT 10.717 20.489 11.609 20.539 ;
		LAYER M4 ;
		RECT 10.717 21.749 11.609 21.799 ;
		LAYER M4 ;
		RECT 10.717 22.505 11.609 22.555 ;
		LAYER M4 ;
		RECT 10.717 23.765 11.609 23.815 ;
		LAYER M4 ;
		RECT 10.717 24.521 11.609 24.571 ;
		LAYER M4 ;
		RECT 10.717 25.781 11.609 25.831 ;
		LAYER M4 ;
		RECT 10.717 26.537 11.609 26.587 ;
		LAYER M4 ;
		RECT 10.717 27.797 11.609 27.847 ;
		LAYER M4 ;
		RECT 10.717 28.553 11.609 28.603 ;
		LAYER M4 ;
		RECT 10.717 29.813 11.609 29.863 ;
		LAYER M4 ;
		RECT 10.717 30.569 11.609 30.619 ;
		LAYER M4 ;
		RECT 10.717 31.829 11.609 31.879 ;
		LAYER M4 ;
		RECT 10.717 32.585 11.609 32.635 ;
		LAYER M4 ;
		RECT 10.717 33.845 11.609 33.895 ;
		LAYER M4 ;
		RECT 10.717 34.601 11.609 34.651 ;
		LAYER M4 ;
		RECT 10.717 35.861 11.609 35.911 ;
		LAYER M4 ;
		RECT 10.717 36.617 11.609 36.667 ;
		LAYER M4 ;
		RECT 10.717 37.877 11.609 37.927 ;
		LAYER M4 ;
		RECT 10.717 38.633 11.609 38.683 ;
		LAYER M4 ;
		RECT 10.717 39.893 11.609 39.943 ;
		LAYER M4 ;
		RECT 10.717 40.649 11.609 40.699 ;
		LAYER M4 ;
		RECT 10.717 41.909 11.609 41.959 ;
		LAYER M4 ;
		RECT 10.717 42.665 11.609 42.715 ;
		LAYER M4 ;
		RECT 10.717 43.925 11.609 43.975 ;
		LAYER M4 ;
		RECT 10.717 44.681 11.609 44.731 ;
		LAYER M4 ;
		RECT 10.717 45.941 11.609 45.991 ;
		LAYER M4 ;
		RECT 10.717 46.697 11.609 46.747 ;
		LAYER M4 ;
		RECT 10.717 47.957 11.609 48.007 ;
		LAYER M4 ;
		RECT 10.717 48.713 11.609 48.763 ;
		LAYER M4 ;
		RECT 10.717 49.973 11.609 50.023 ;
		LAYER M4 ;
		RECT 10.717 50.729 11.609 50.779 ;
		LAYER M4 ;
		RECT 10.717 51.989 11.609 52.039 ;
		LAYER M4 ;
		RECT 10.717 52.745 11.609 52.795 ;
		LAYER M4 ;
		RECT 10.717 54.005 11.609 54.055 ;
		LAYER M4 ;
		RECT 10.717 54.761 11.609 54.811 ;
		LAYER M4 ;
		RECT 10.717 56.021 11.609 56.071 ;
		LAYER M4 ;
		RECT 10.717 56.777 11.609 56.827 ;
		LAYER M4 ;
		RECT 10.717 58.037 11.609 58.087 ;
		LAYER M4 ;
		RECT 10.717 58.793 11.609 58.843 ;
		LAYER M4 ;
		RECT 10.717 60.053 11.609 60.103 ;
		LAYER M4 ;
		RECT 10.717 60.809 11.609 60.859 ;
		LAYER M4 ;
		RECT 10.717 62.069 11.609 62.119 ;
		LAYER M4 ;
		RECT 10.717 62.825 11.609 62.875 ;
		LAYER M4 ;
		RECT 10.717 64.085 11.609 64.135 ;
		LAYER M4 ;
		RECT 10.717 64.841 11.609 64.891 ;
		LAYER M4 ;
		RECT 10.717 66.101 11.609 66.151 ;
		LAYER M4 ;
		RECT 10.717 66.857 11.609 66.907 ;
		LAYER M4 ;
		RECT 10.717 68.117 11.609 68.167 ;
		LAYER M4 ;
		RECT 10.717 68.873 11.609 68.923 ;
		LAYER M4 ;
		RECT 10.717 70.133 11.609 70.183 ;
		LAYER M4 ;
		RECT 10.717 70.889 11.609 70.939 ;
		LAYER M4 ;
		RECT 10.717 72.149 11.609 72.199 ;
		LAYER M4 ;
		RECT 10.717 72.905 11.609 72.955 ;
		LAYER M4 ;
		RECT 10.717 74.165 11.609 74.215 ;
		LAYER M4 ;
		RECT 10.717 74.921 11.609 74.971 ;
		LAYER M4 ;
		RECT 10.717 76.181 11.609 76.231 ;
		LAYER M4 ;
		RECT 10.717 76.937 11.609 76.987 ;
		LAYER M4 ;
		RECT 10.717 78.197 11.609 78.247 ;
		LAYER M4 ;
		RECT 10.717 78.953 11.609 79.003 ;
		LAYER M4 ;
		RECT 10.717 80.213 11.609 80.263 ;
		LAYER M4 ;
		RECT 10.717 80.969 11.609 81.019 ;
		LAYER M4 ;
		RECT 10.717 82.229 11.609 82.279 ;
		LAYER M4 ;
		RECT 10.717 82.985 11.609 83.035 ;
		LAYER M4 ;
		RECT 10.717 84.245 11.609 84.295 ;
		LAYER M4 ;
		RECT 10.717 85.001 11.609 85.051 ;
		LAYER M4 ;
		RECT 10.717 86.261 11.609 86.311 ;
		LAYER M4 ;
		RECT 10.717 87.017 11.609 87.067 ;
		LAYER M4 ;
		RECT 10.717 88.277 11.609 88.327 ;
		LAYER M4 ;
		RECT 10.717 89.033 11.609 89.083 ;
		LAYER M4 ;
		RECT 10.717 90.293 11.609 90.343 ;
		LAYER M4 ;
		RECT 10.717 91.049 11.609 91.099 ;
		LAYER M4 ;
		RECT 10.717 92.309 11.609 92.359 ;
		LAYER M4 ;
		RECT 10.717 93.065 11.609 93.115 ;
		LAYER M4 ;
		RECT 10.717 94.325 11.609 94.375 ;
		LAYER M4 ;
		RECT 10.717 95.081 11.609 95.131 ;
		LAYER M4 ;
		RECT 10.717 96.341 11.609 96.391 ;
		LAYER M4 ;
		RECT 10.717 97.097 11.609 97.147 ;
		LAYER M4 ;
		RECT 10.717 98.357 11.609 98.407 ;
		LAYER M4 ;
		RECT 10.717 99.113 11.609 99.163 ;
		LAYER M4 ;
		RECT 10.717 100.373 11.609 100.423 ;
		LAYER M4 ;
		RECT 10.717 101.129 11.609 101.179 ;
		LAYER M4 ;
		RECT 10.717 102.389 11.609 102.439 ;
		LAYER M4 ;
		RECT 10.717 103.145 11.609 103.195 ;
		LAYER M4 ;
		RECT 10.717 104.405 11.609 104.455 ;
		LAYER M4 ;
		RECT 10.717 105.161 11.609 105.211 ;
		LAYER M4 ;
		RECT 10.717 106.421 11.609 106.471 ;
		LAYER M4 ;
		RECT 10.717 107.177 11.609 107.227 ;
		LAYER M4 ;
		RECT 10.717 108.437 11.609 108.487 ;
		LAYER M4 ;
		RECT 10.717 109.193 11.609 109.243 ;
		LAYER M4 ;
		RECT 10.717 110.453 11.609 110.503 ;
		LAYER M4 ;
		RECT 10.717 111.209 11.609 111.259 ;
		LAYER M4 ;
		RECT 10.717 112.469 11.609 112.519 ;
		LAYER M4 ;
		RECT 10.717 113.225 11.609 113.275 ;
		LAYER M4 ;
		RECT 10.717 114.485 11.609 114.535 ;
		LAYER M4 ;
		RECT 10.717 115.241 11.609 115.291 ;
		LAYER M4 ;
		RECT 10.717 116.501 11.609 116.551 ;
		LAYER M4 ;
		RECT 10.717 117.257 11.609 117.307 ;
		LAYER M4 ;
		RECT 10.717 118.517 11.609 118.567 ;
		LAYER M4 ;
		RECT 10.717 119.273 11.609 119.323 ;
		LAYER M4 ;
		RECT 10.717 120.533 11.609 120.583 ;
		LAYER M4 ;
		RECT 10.717 121.289 11.609 121.339 ;
		LAYER M4 ;
		RECT 10.717 122.549 11.609 122.599 ;
		LAYER M4 ;
		RECT 10.717 123.305 11.609 123.355 ;
		LAYER M4 ;
		RECT 10.717 124.565 11.609 124.615 ;
		LAYER M4 ;
		RECT 10.717 125.321 11.609 125.371 ;
		LAYER M4 ;
		RECT 10.717 126.581 11.609 126.631 ;
		LAYER M4 ;
		RECT 10.717 127.337 11.609 127.387 ;
		LAYER M4 ;
		RECT 10.717 128.597 11.609 128.647 ;
		LAYER M4 ;
		RECT 10.717 129.353 11.609 129.403 ;
		LAYER M4 ;
		RECT 10.717 143.477 11.609 143.527 ;
		LAYER M4 ;
		RECT 10.717 144.233 11.609 144.283 ;
		LAYER M4 ;
		RECT 10.717 145.493 11.609 145.543 ;
		LAYER M4 ;
		RECT 10.717 146.249 11.609 146.299 ;
		LAYER M4 ;
		RECT 10.717 147.509 11.609 147.559 ;
		LAYER M4 ;
		RECT 10.717 148.265 11.609 148.315 ;
		LAYER M4 ;
		RECT 10.717 149.525 11.609 149.575 ;
		LAYER M4 ;
		RECT 10.717 150.281 11.609 150.331 ;
		LAYER M4 ;
		RECT 10.717 151.541 11.609 151.591 ;
		LAYER M4 ;
		RECT 10.717 152.297 11.609 152.347 ;
		LAYER M4 ;
		RECT 10.717 153.557 11.609 153.607 ;
		LAYER M4 ;
		RECT 10.717 154.313 11.609 154.363 ;
		LAYER M4 ;
		RECT 10.717 155.573 11.609 155.623 ;
		LAYER M4 ;
		RECT 10.717 156.329 11.609 156.379 ;
		LAYER M4 ;
		RECT 10.717 157.589 11.609 157.639 ;
		LAYER M4 ;
		RECT 10.717 158.345 11.609 158.395 ;
		LAYER M4 ;
		RECT 10.717 159.605 11.609 159.655 ;
		LAYER M4 ;
		RECT 10.717 160.361 11.609 160.411 ;
		LAYER M4 ;
		RECT 10.717 161.621 11.609 161.671 ;
		LAYER M4 ;
		RECT 10.717 162.377 11.609 162.427 ;
		LAYER M4 ;
		RECT 10.717 163.637 11.609 163.687 ;
		LAYER M4 ;
		RECT 10.717 164.393 11.609 164.443 ;
		LAYER M4 ;
		RECT 10.717 165.653 11.609 165.703 ;
		LAYER M4 ;
		RECT 10.717 166.409 11.609 166.459 ;
		LAYER M4 ;
		RECT 10.717 167.669 11.609 167.719 ;
		LAYER M4 ;
		RECT 10.717 168.425 11.609 168.475 ;
		LAYER M4 ;
		RECT 10.717 169.685 11.609 169.735 ;
		LAYER M4 ;
		RECT 10.717 170.441 11.609 170.491 ;
		LAYER M4 ;
		RECT 10.717 171.701 11.609 171.751 ;
		LAYER M4 ;
		RECT 10.717 172.457 11.609 172.507 ;
		LAYER M4 ;
		RECT 10.717 173.717 11.609 173.767 ;
		LAYER M4 ;
		RECT 10.717 174.473 11.609 174.523 ;
		LAYER M4 ;
		RECT 10.717 175.733 11.609 175.783 ;
		LAYER M4 ;
		RECT 10.717 176.489 11.609 176.539 ;
		LAYER M4 ;
		RECT 10.717 177.749 11.609 177.799 ;
		LAYER M4 ;
		RECT 10.717 178.505 11.609 178.555 ;
		LAYER M4 ;
		RECT 10.717 179.765 11.609 179.815 ;
		LAYER M4 ;
		RECT 10.717 180.521 11.609 180.571 ;
		LAYER M4 ;
		RECT 10.717 181.781 11.609 181.831 ;
		LAYER M4 ;
		RECT 10.717 182.537 11.609 182.587 ;
		LAYER M4 ;
		RECT 10.717 183.797 11.609 183.847 ;
		LAYER M4 ;
		RECT 10.717 184.553 11.609 184.603 ;
		LAYER M4 ;
		RECT 10.717 185.813 11.609 185.863 ;
		LAYER M4 ;
		RECT 10.717 186.569 11.609 186.619 ;
		LAYER M4 ;
		RECT 10.717 187.829 11.609 187.879 ;
		LAYER M4 ;
		RECT 10.717 188.585 11.609 188.635 ;
		LAYER M4 ;
		RECT 10.717 189.845 11.609 189.895 ;
		LAYER M4 ;
		RECT 10.717 190.601 11.609 190.651 ;
		LAYER M4 ;
		RECT 10.717 191.861 11.609 191.911 ;
		LAYER M4 ;
		RECT 10.717 192.617 11.609 192.667 ;
		LAYER M4 ;
		RECT 10.717 193.877 11.609 193.927 ;
		LAYER M4 ;
		RECT 10.717 194.633 11.609 194.683 ;
		LAYER M4 ;
		RECT 10.717 195.893 11.609 195.943 ;
		LAYER M4 ;
		RECT 10.717 196.649 11.609 196.699 ;
		LAYER M4 ;
		RECT 10.717 197.909 11.609 197.959 ;
		LAYER M4 ;
		RECT 10.717 198.665 11.609 198.715 ;
		LAYER M4 ;
		RECT 10.717 199.925 11.609 199.975 ;
		LAYER M4 ;
		RECT 10.717 200.681 11.609 200.731 ;
		LAYER M4 ;
		RECT 10.717 201.941 11.609 201.991 ;
		LAYER M4 ;
		RECT 10.717 202.697 11.609 202.747 ;
		LAYER M4 ;
		RECT 10.717 203.957 11.609 204.007 ;
		LAYER M4 ;
		RECT 10.717 204.713 11.609 204.763 ;
		LAYER M4 ;
		RECT 10.717 205.973 11.609 206.023 ;
		LAYER M4 ;
		RECT 10.717 206.729 11.609 206.779 ;
		LAYER M4 ;
		RECT 10.717 207.989 11.609 208.039 ;
		LAYER M4 ;
		RECT 10.717 208.745 11.609 208.795 ;
		LAYER M4 ;
		RECT 10.717 210.005 11.609 210.055 ;
		LAYER M4 ;
		RECT 10.717 210.761 11.609 210.811 ;
		LAYER M4 ;
		RECT 10.717 212.021 11.609 212.071 ;
		LAYER M4 ;
		RECT 10.717 212.777 11.609 212.827 ;
		LAYER M4 ;
		RECT 10.717 214.037 11.609 214.087 ;
		LAYER M4 ;
		RECT 10.717 214.793 11.609 214.843 ;
		LAYER M4 ;
		RECT 10.717 216.053 11.609 216.103 ;
		LAYER M4 ;
		RECT 10.717 216.809 11.609 216.859 ;
		LAYER M4 ;
		RECT 10.717 218.069 11.609 218.119 ;
		LAYER M4 ;
		RECT 10.717 218.825 11.609 218.875 ;
		LAYER M4 ;
		RECT 10.717 220.085 11.609 220.135 ;
		LAYER M4 ;
		RECT 10.717 220.841 11.609 220.891 ;
		LAYER M4 ;
		RECT 10.717 222.101 11.609 222.151 ;
		LAYER M4 ;
		RECT 10.717 222.857 11.609 222.907 ;
		LAYER M4 ;
		RECT 10.717 224.117 11.609 224.167 ;
		LAYER M4 ;
		RECT 10.717 224.873 11.609 224.923 ;
		LAYER M4 ;
		RECT 10.717 226.133 11.609 226.183 ;
		LAYER M4 ;
		RECT 10.717 226.889 11.609 226.939 ;
		LAYER M4 ;
		RECT 10.717 228.149 11.609 228.199 ;
		LAYER M4 ;
		RECT 10.717 228.905 11.609 228.955 ;
		LAYER M4 ;
		RECT 10.717 230.165 11.609 230.215 ;
		LAYER M4 ;
		RECT 10.717 230.921 11.609 230.971 ;
		LAYER M4 ;
		RECT 10.717 232.181 11.609 232.231 ;
		LAYER M4 ;
		RECT 10.717 232.937 11.609 232.987 ;
		LAYER M4 ;
		RECT 10.717 234.197 11.609 234.247 ;
		LAYER M4 ;
		RECT 10.717 234.953 11.609 235.003 ;
		LAYER M4 ;
		RECT 10.717 236.213 11.609 236.263 ;
		LAYER M4 ;
		RECT 10.717 236.969 11.609 237.019 ;
		LAYER M4 ;
		RECT 10.717 238.229 11.609 238.279 ;
		LAYER M4 ;
		RECT 10.717 238.985 11.609 239.035 ;
		LAYER M4 ;
		RECT 10.717 240.245 11.609 240.295 ;
		LAYER M4 ;
		RECT 10.717 241.001 11.609 241.051 ;
		LAYER M4 ;
		RECT 10.717 242.261 11.609 242.311 ;
		LAYER M4 ;
		RECT 10.717 243.017 11.609 243.067 ;
		LAYER M4 ;
		RECT 10.717 244.277 11.609 244.327 ;
		LAYER M4 ;
		RECT 10.717 245.033 11.609 245.083 ;
		LAYER M4 ;
		RECT 10.717 246.293 11.609 246.343 ;
		LAYER M4 ;
		RECT 10.717 247.049 11.609 247.099 ;
		LAYER M4 ;
		RECT 10.717 248.309 11.609 248.359 ;
		LAYER M4 ;
		RECT 10.717 249.065 11.609 249.115 ;
		LAYER M4 ;
		RECT 10.717 250.325 11.609 250.375 ;
		LAYER M4 ;
		RECT 10.717 251.081 11.609 251.131 ;
		LAYER M4 ;
		RECT 10.717 252.341 11.609 252.391 ;
		LAYER M4 ;
		RECT 10.717 253.097 11.609 253.147 ;
		LAYER M4 ;
		RECT 10.717 254.357 11.609 254.407 ;
		LAYER M4 ;
		RECT 10.717 255.113 11.609 255.163 ;
		LAYER M4 ;
		RECT 10.717 256.373 11.609 256.423 ;
		LAYER M4 ;
		RECT 10.717 257.129 11.609 257.179 ;
		LAYER M4 ;
		RECT 10.717 258.389 11.609 258.439 ;
		LAYER M4 ;
		RECT 10.717 259.145 11.609 259.195 ;
		LAYER M4 ;
		RECT 10.717 260.405 11.609 260.455 ;
		LAYER M4 ;
		RECT 10.717 261.161 11.609 261.211 ;
		LAYER M4 ;
		RECT 10.717 262.421 11.609 262.471 ;
		LAYER M4 ;
		RECT 10.717 263.177 11.609 263.227 ;
		LAYER M4 ;
		RECT 10.717 264.437 11.609 264.487 ;
		LAYER M4 ;
		RECT 10.717 265.193 11.609 265.243 ;
		LAYER M4 ;
		RECT 10.717 266.453 11.609 266.503 ;
		LAYER M4 ;
		RECT 10.717 267.209 11.609 267.259 ;
		LAYER M4 ;
		RECT 10.717 268.469 11.609 268.519 ;
		LAYER M4 ;
		RECT 10.717 269.225 11.609 269.275 ;
		LAYER M4 ;
		RECT 10.717 270.485 11.609 270.535 ;
		LAYER M4 ;
		RECT 10.717 271.241 11.609 271.291 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 17.375 272.880 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 17.375 272.880 ;
	END
END TS1N16FFCLLSVTA64X128M4SW

END LIBRARY
