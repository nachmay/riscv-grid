**** Created by MC2: Version 2013.12.00.f on 2025/06/18, 13:11:27 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  TS16FF2PRF
* Top Cell Name: all_leafcells
* View Name:     schematic
* Netlisted on:  Sep 30 16:22:09 2015
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM


*.PIN vss

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_svt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nand2_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_svt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_inv_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_svt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nor2_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WCTD VDD VDDI VSS TSMC_1 TSMC_2 TSMC_3 TSMC_4 
XI76 TSMC_5 TSMC_6 VSS VSS VDDI VDD TSMC_3 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI79 TSMC_7 TSMC_8 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI66 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_2 TSMC_11 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_7 TSMC_12 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_14 TSMC_7 VSS VSS VDDI VDD TSMC_6 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_1 TSMC_15 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_9 TSMC_16 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_17 TSMC_11 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_16 TSMC_15 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI145 VSS VSS TSMC_4 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_18 TSMC_5 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_5 TSMC_19 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_5 TSMC_20 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI143 VSS VSS TSMC_21 TSMC_22 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI159 VSS VSS TSMC_13 TSMC_23 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_22 TSMC_17 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_24 TSMC_25 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI89 VSS VSS TSMC_10 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI160 VSS VSS TSMC_13 TSMC_24 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI144 VSS VSS TSMC_25 TSMC_21 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI64 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW8U20_nor2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WRTRKEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WRTRKEN TSMC_1 VDD VDDI VSS TSMC_2 TSMC_3 TSMC_4 
XI19<0> TSMC_2 TSMC_5 VSS VSS VDDI VDD TSMC_1 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI19<1> TSMC_2 TSMC_5 VSS VSS VDDI VDD TSMC_1 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI14 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_5 
+ S6ALLSVTFW8U20_nor2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_W1TRKWR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_W1TRKWR TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS TSMC_4 
+ TSMC_5 
XXwctd VDD VDDI VSS TSMC_1 TSMC_2 TSMC_6 TSMC_4 S6ALLSVTFW8U20_RF_WCTD 
XXrdtrken TSMC_3 VDD VDDI VSS TSMC_6 TSMC_4 TSMC_5 
+ S6ALLSVTFW8U20_RF_WRTRKEN 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WREFMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WREFMUX TSMC_1 VDD VDDI VSS TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
MM10 TSMC_7 TSMC_1 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_4 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_4 TSMC_6 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM13 TSMC_8 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_3 TSMC_6 TSMC_9 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM12 TSMC_9 TSMC_1 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_3 TSMC_5 TSMC_4 VDD pch_svt_mac l=0.020u nfin=3 m=2 
MM9 TSMC_3 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM8 TSMC_4 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM0 TSMC_3 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_1 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_3 TSMC_10 TSMC_2 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM5 TSMC_4 TSMC_11 TSMC_2 VSS nch_svt_mac l=0.020u nfin=6 m=2 
XI21 TSMC_6 TSMC_7 TSMC_2 VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI19 TSMC_6 TSMC_1 TSMC_2 VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKGIOWR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TRKGIOWR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 
XXwrst TSMC_15 TSMC_16 TSMC_20 VDD VDDI VSS TSMC_17 TSMC_29 
+ S6ALLSVTFW8U20_RF_W1TRKWR 
XXwrefmux TSMC_11 VDD VDDI VSS VSS TSMC_12 TSMC_14 TSMC_30 TSMC_29 
+ S6ALLSVTFW8U20_RF_WREFMUX 
XI21 VSS VSS TSMC_19 TSMC_29 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_29 TSMC_30 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 p_nfin=7 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WMUX TSMC_1 TSMC_2 VDD VDDI VSS TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM0 TSMC_4 TSMC_8 TSMC_3 VSS nch_lvt_mac l=0.020u nfin=6 m=2 
MM2 TSMC_5 TSMC_9 TSMC_3 VSS nch_lvt_mac l=0.020u nfin=6 m=2 
MM13 TSMC_10 TSMC_1 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_4 TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_4 TSMC_11 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_5 TSMC_11 TSMC_10 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM9 TSMC_4 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM4 TSMC_5 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=6 m=2 
MM10 TSMC_4 TSMC_6 TSMC_5 VDD pch_svt_mac l=0.020u nfin=3 m=2 
MM6 TSMC_5 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM12 TSMC_12 TSMC_2 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI23 VSS VSS TSMC_7 TSMC_11 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI14 TSMC_11 TSMC_2 TSMC_3 VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI15 TSMC_11 TSMC_1 TSMC_3 VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRI_W3L2M1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TRI_W3L2M1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM4 TSMC_9 TSMC_7 TSMC_4 TSMC_5 pch_svt_mac l=0.020u nfin=3 m=1 
MM5 TSMC_8 TSMC_1 TSMC_9 TSMC_5 pch_svt_mac l=0.020u nfin=3 m=1 
MM6 TSMC_10 TSMC_6 TSMC_2 TSMC_3 nch_svt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_8 TSMC_1 TSMC_10 TSMC_3 nch_svt_mac l=0.020u nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRI_W2L2M1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TRI_W2L2M1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
MM4 TSMC_9 TSMC_7 TSMC_4 TSMC_5 pch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_8 TSMC_1 TSMC_9 TSMC_5 pch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_10 TSMC_6 TSMC_2 TSMC_3 nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_8 TSMC_1 TSMC_10 TSMC_3 nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DIN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_DIN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD 
+ VDDI VSS TSMC_7 
XI16 TSMC_8 VSS VSS VDDI VDD TSMC_4 TSMC_5 TSMC_9 
+ S6ALLSVTFW8U20_RF_TRI_W3L2M1 
XI90 TSMC_10 VSS VSS VDDI VDD TSMC_4 TSMC_5 TSMC_11 
+ S6ALLSVTFW8U20_RF_TRI_W3L2M1 
XI15 TSMC_12 TSMC_13 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_12 TSMC_14 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI63 VSS VSS TSMC_15 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI59 VSS VSS TSMC_16 TSMC_14 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI61 VSS VSS TSMC_7 TSMC_17 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI83 VSS VSS TSMC_9 TSMC_3 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI92 VSS VSS TSMC_11 TSMC_2 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI99 VSS VSS TSMC_1 TSMC_16 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI62 VSS VSS TSMC_17 TSMC_15 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI60 VSS VSS TSMC_14 TSMC_13 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI94 TSMC_2 VSS VSS VDDI VDD TSMC_5 TSMC_4 TSMC_11 
+ S6ALLSVTFW8U20_RF_TRI_W2L2M1 
XI17 TSMC_3 VSS VSS VDDI VDD TSMC_5 TSMC_4 TSMC_9 
+ S6ALLSVTFW8U20_RF_TRI_W2L2M1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    TRI_M2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_TRI_M2 TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS TSMC_4 
MM4 TSMC_5 TSMC_1 VDDI VDD pch_lvt_mac l=0.020u nfin=4 m=1 
MM5 TSMC_4 TSMC_3 TSMC_5 VDD pch_lvt_mac l=0.020u nfin=4 m=1 
MM6 TSMC_6 TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=4 m=1 
MM3 TSMC_4 TSMC_2 TSMC_6 VSS nch_svt_mac l=0.020u nfin=4 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RMUX
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RMUX TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI VSS 
XI9 TSMC_1 TSMC_5 TSMC_4 VDD VDDI VSS TSMC_2 S6ALLSVTFW8U20_TRI_M2 
MM2 TSMC_1 TSMC_6 TSMC_7 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_7 TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_1 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=4 m=3 
MM5 TSMC_8 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_1 TSMC_6 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI1 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DOLATCH
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_DOLATCH TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD 
+ VDDI VSS TSMC_7 TSMC_8 
MM2 TSMC_3 TSMC_4 VDD VDD pch_svt_mac l=0.020u nfin=3 m=1 
XI3 VSS VSS TSMC_3 TSMC_1 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI7 TSMC_2 VSS VSS VDDI VDD TSMC_5 TSMC_6 TSMC_3 
+ S6ALLSVTFW8U20_RF_TRI_W2L2M1 
XI5 TSMC_3 VSS VSS VDDI VDD TSMC_7 TSMC_8 TSMC_2 
+ S6ALLSVTFW8U20_RF_TRI_W2L2M1 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_svt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nand3_svt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RLCTRL_DK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RLCTRL_DK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 VDD VDDI VSS TSMC_27 
MM12 TSMC_28 TSMC_29 TSMC_30 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM11 TSMC_30 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM7 TSMC_32 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM6 TSMC_33 TSMC_34 TSMC_32 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM5 TSMC_33 TSMC_35 TSMC_32 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM1 TSMC_36 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=8 m=16 
MM0 TSMC_36 TSMC_31 VSS VSS nch_ulvt_mac l=0.020u nfin=8 m=16 
MM8 TSMC_28 TSMC_35 TSMC_30 VSS nch_ulvt_mac l=0.020u nfin=2 m=3 
MM13 TSMC_28 TSMC_31 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM4 TSMC_33 TSMC_31 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM3 TSMC_33 TSMC_35 TSMC_37 VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM2 TSMC_37 TSMC_34 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM10 TSMC_38 TSMC_29 VDD VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
MM9 TSMC_28 TSMC_35 TSMC_38 VDD pch_ulvt_mac l=0.020u nfin=3 m=3 
XI96 TSMC_36 VSS TSMC_39 TSMC_18 VDD VDD 
+ S6ALLSVTFW8U20_inv_ulvt_mac_pcell n_totalM=16 n_nfin=6 n_l=0.020u p_totalM=16 
+ p_nfin=6 p_l=0.020u 
XI100 VSS VSS TSMC_1 TSMC_40 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=5 p_l=0.020u 
XI107 VSS VSS TSMC_41 TSMC_5 VDD VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI91 VSS VSS TSMC_33 TSMC_42 VDD VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=5 n_nfin=7 n_l=0.020u p_totalM=5 p_nfin=6 p_l=0.020u 
XI92 TSMC_36 VSS TSMC_42 TSMC_19 VDD VDD 
+ S6ALLSVTFW8U20_inv_ulvt_mac_pcell n_totalM=16 n_nfin=6 n_l=0.020u p_totalM=16 
+ p_nfin=6 p_l=0.020u 
XI106 VSS VSS TSMC_4 TSMC_41 VDD VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI98 VSS VSS TSMC_35 TSMC_23 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=14 n_nfin=5 n_l=0.020u p_totalM=14 p_nfin=5 p_l=0.020u 
XI101 VSS VSS TSMC_40 TSMC_11 VDDI VDD 
+ S6ALLSVTFW8U20_inv_ulvt_mac_pcell n_totalM=10 n_nfin=7 n_l=0.020u p_totalM=10 
+ p_nfin=8 p_l=0.020u 
XI93_Lg16 TSMC_21 TSMC_22 TSMC_27 VSS VSS VDD VDD TSMC_35 
+ S6ALLSVTFW8U20_nand3_ulvt_mac_pcell n_totalM=4 n_nfin=7 n_l=0.020u p_totalM=4 
+ p_nfin=2 p_l=0.020u 
XI95 TSMC_25 TSMC_26 VSS VSS VDDI VDD TSMC_34 
+ S6ALLSVTFW8U20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI103 TSMC_28 TSMC_24 VSS VSS VDD VDD TSMC_39 
+ S6ALLSVTFW8U20_nor2_ulvt_mac_pcell n_totalM=6 n_nfin=6 n_l=0.020u p_totalM=6 
+ p_nfin=7 p_l=0.020u 
XI102 TSMC_4 TSMC_4 VSS VSS VDD VDD TSMC_31 
+ S6ALLSVTFW8U20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI99 TSMC_2 TSMC_3 VSS VSS VDDI VDD TSMC_29 
+ S6ALLSVTFW8U20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WLCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WLCTRL VDD VDDI VSS TSMC_1 TSMC_2 TSMC_3 TSMC_4 
XI27 TSMC_1 TSMC_2 TSMC_4 VSS VSS VDD VDD TSMC_5 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=4 n_nfin=7 n_l=0.020u p_totalM=4 
+ p_nfin=2 p_l=0.020u 
XI28 VSS VSS TSMC_5 TSMC_3 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=14 n_nfin=5 n_l=0.020u p_totalM=14 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LCTRL_DK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_LCTRL_DK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
MM6 TSMC_71 TSMC_46 VDD VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM4 VDDI TSMC_46 VDDI VDD pch_ulvt_mac l=0.020u nfin=8 m=2 
MM5 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=12 m=16 
MM1 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=5 m=16 
MM0 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=9 m=32 
MM2 VDDI TSMC_72 VDD VDD pch_svt_mac l=0.020u nfin=10 m=16 
XXrlctrl TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_17 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_25 TSMC_27 TSMC_28 TSMC_45 TSMC_48 TSMC_49 VDD 
+ VDDI VSS TSMC_69 S6ALLSVTFW8U20_RF_RLCTRL_DK 
XXwlctrl VDD VDDI VSS TSMC_50 TSMC_51 TSMC_52 TSMC_70 
+ S6ALLSVTFW8U20_RF_WLCTRL 
XI51 VSS VSS TSMC_73 TSMC_72 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI52 TSMC_24 TSMC_4 VSS VSS VDD VDD TSMC_73 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
MM3 VSS TSMC_46 VSS VSS nch_ulvt_mac l=0.020u nfin=7 m=2 
MM7 TSMC_46 TSMC_71 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_LCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
XI152 TSMC_15 TSMC_24 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=2 n_nfin=12 n_l=0.020u p_totalM=2 
+ p_nfin=12 p_l=0.020u 
XI49<1> VSS VSS TSMC_18 TSMC_12 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI49<0> VSS VSS TSMC_19 TSMC_13 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
Xlctrl TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 VDD VDDI VSS 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ S6ALLSVTFW8U20_RF_LCTRL_DK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_XDECCAP
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_XDECCAP TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 
MM0_LVT TSMC_12 TSMC_6 VSS VSS nch_lvt_mac l=0.020u nfin=5 m=1 
MM196_LVT TSMC_13 TSMC_12 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM197_LVT TSMC_14 TSMC_12 TSMC_13 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM194_LVT TSMC_12 TSMC_15 VSS VSS nch_lvt_mac l=0.020u nfin=5 m=1 
MM4 TSMC_10 TSMC_16 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MMWLDRPCHWTK TSMC_10 TSMC_16 VDDI VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM195_LVT TSMC_14 TSMC_12 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=2 
MM198_LVT TSMC_17 TSMC_15 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM193_LVT TSMC_12 TSMC_6 TSMC_17 VDD pch_lvt_mac l=0.020u nfin=2 m=1 
XI78 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=6 n_l=0.020u p_totalM=2 p_nfin=6 p_l=0.020u 
XI75 VSS VSS TSMC_9 TSMC_18 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI79 VSS VSS TSMC_3 TSMC_4 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI72_LVT VSS VSS TSMC_11 TSMC_15 VDDI VDD 
+ S6ALLSVTFW8U20_inv_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI73_LVT VSS VSS TSMC_14 TSMC_19 VDDI VDD 
+ S6ALLSVTFW8U20_inv_lvt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI77 VSS VSS TSMC_2 TSMC_20 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI76 VSS VSS TSMC_18 TSMC_21 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=2 p_l=0.020u 
XI81_LVT TSMC_10 TSMC_19 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=8 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
XI82 TSMC_20 TSMC_21 VSS VSS VDD VDD TSMC_16 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=12 n_l=0.020u p_totalM=1 
+ p_nfin=10 p_l=0.020u 
XI80_LVT TSMC_10 TSMC_19 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=6 n_l=0.020u p_totalM=1 
+ p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TRKCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 VDD VDDI VSS TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 
MM4 TSMC_37 TSMC_56 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
XI76 VSS VSS TSMC_57 TSMC_58 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI75 VSS VSS TSMC_12 TSMC_57 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI78 TSMC_13 TSMC_14 VSS VSS VDD VDD TSMC_56 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=12 n_l=0.020u p_totalM=1 
+ p_nfin=6 p_l=0.020u 
XI79 TSMC_58 TSMC_14 VSS VSS VDDI VDD TSMC_59 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=7 p_l=0.020u 
MMWLDRPCHRTK TSMC_37 TSMC_56 VDDI VDD pch_svt_mac l=0.020u nfin=11 m=4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DOUTM1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_DOUTM1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS TSMC_11 TSMC_12 
XXqltch TSMC_5 TSMC_1 TSMC_13 TSMC_4 TSMC_6 TSMC_7 VDD VDDI VSS TSMC_11 TSMC_12 
+ S6ALLSVTFW8U20_RF_DOLATCH 
XXrmux<0> TSMC_2 TSMC_13 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS 
+ S6ALLSVTFW8U20_RF_RMUX 
XI26 VSS VSS TSMC_3 TSMC_4 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DINM1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_DINM1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
XXdltch TSMC_1 TSMC_11 TSMC_12 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS TSMC_8 
+ S6ALLSVTFW8U20_RF_DIN 
XXwmux<0> TSMC_11 TSMC_12 VDD VDDI VSS TSMC_5 TSMC_6 TSMC_7 TSMC_9 TSMC_10 
+ S6ALLSVTFW8U20_RF_WMUX 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_GIOM1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_GIOM1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 VDD VDDI VSS 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 
XXdout TSMC_2 TSMC_3 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 VDD VDDI VSS TSMC_16 TSMC_17 S6ALLSVTFW8U20_RF_DOUTM1 
XXdin TSMC_1 TSMC_4 TSMC_5 TSMC_14 VDD VDDI VSS TSMC_15 TSMC_18 TSMC_19 TSMC_20 
+ TSMC_21 TSMC_26 S6ALLSVTFW8U20_RF_DINM1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_GIOM1X2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_GIOM1X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 
XXgio1 TSMC_1 TSMC_3 TSMC_5 TSMC_30 TSMC_31 TSMC_7 TSMC_32 TSMC_8 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_11 VDD VDDI VSS TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_18 TSMC_20 TSMC_38 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 TSMC_28 S6ALLSVTFW8U20_RF_GIOM1 
XXgio0 TSMC_2 TSMC_4 TSMC_6 TSMC_30 TSMC_31 TSMC_7 TSMC_32 TSMC_9 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_11 VDD VDDI VSS TSMC_12 TSMC_14 
+ TSMC_15 TSMC_17 TSMC_19 TSMC_21 TSMC_38 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 TSMC_29 S6ALLSVTFW8U20_RF_GIOM1 
XI25 VSS VSS TSMC_34 TSMC_33 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI32 VSS VSS TSMC_34 TSMC_39 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI26 VSS VSS TSMC_40 TSMC_37 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI11 VSS VSS TSMC_30 TSMC_31 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_22 TSMC_30 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI7 VSS VSS TSMC_41 TSMC_38 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 p_nfin=6 p_l=0.020u 
XI5 VSS VSS TSMC_23 TSMC_41 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI23 VSS VSS TSMC_37 TSMC_36 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI28 VSS VSS TSMC_39 TSMC_35 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI34 TSMC_14 TSMC_10 VSS VSS VDD VDD TSMC_40 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI20 TSMC_40 TSMC_32 VSS VSS VDD VDD TSMC_34 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WXDEC TSMC_1 TSMC_2 TSMC_3 VDD VDDI TSMC_4 VSS TSMC_5 
+ TSMC_6 
MM3 TSMC_1 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM2 TSMC_7 TSMC_8 TSMC_1 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM4 TSMC_5 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MMWLDRPCH TSMC_5 TSMC_7 TSMC_4 VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MM0 TSMC_7 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
XI58<1> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI58<0> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDECX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WXDECX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD 
+ VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XI64<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XIXDEC<3> TSMC_16 TSMC_2 TSMC_3 VDD VDDI TSMC_7 VSS TSMC_8 TSMC_15 
+ S6ALLSVTFW8U20_RF_WXDEC 
XIXDEC<1> TSMC_16 TSMC_2 TSMC_5 VDD VDDI TSMC_7 VSS TSMC_10 TSMC_15 
+ S6ALLSVTFW8U20_RF_WXDEC 
XIXDEC<0> TSMC_17 TSMC_1 TSMC_6 VDD VDDI TSMC_7 VSS TSMC_11 TSMC_14 
+ S6ALLSVTFW8U20_RF_WXDEC 
XIXDEC<2> TSMC_17 TSMC_1 TSMC_4 VDD VDDI TSMC_7 VSS TSMC_9 TSMC_14 
+ S6ALLSVTFW8U20_RF_WXDEC 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WXDECX4_LR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WXDECX4_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD VDDI TSMC_7 VSS 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ S6ALLSVTFW8U20_RF_WXDECX4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RXDEC TSMC_1 TSMC_2 TSMC_3 VDD VDDI TSMC_4 VSS TSMC_5 
+ TSMC_6 
MM1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MMWLDRPCH TSMC_5 TSMC_7 TSMC_4 VDD pch_svt_mac l=0.020u nfin=11 m=4 
MM0 TSMC_7 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=5 m=2 
MM4 TSMC_5 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=10 m=4 
MM2 TSMC_7 TSMC_8 TSMC_1 VSS nch_svt_mac l=0.020u nfin=6 m=2 
MM3 TSMC_1 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=6 m=2 
XI58<1> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI58<0> TSMC_6 TSMC_3 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDECX4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RXDECX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD 
+ VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC<1> TSMC_14 TSMC_2 TSMC_5 VDD VDDI TSMC_7 VSS TSMC_10 TSMC_15 
+ S6ALLSVTFW8U20_RF_RXDEC 
XIXDEC<3> TSMC_14 TSMC_2 TSMC_3 VDD VDDI TSMC_7 VSS TSMC_8 TSMC_15 
+ S6ALLSVTFW8U20_RF_RXDEC 
XIXDEC<2> TSMC_16 TSMC_1 TSMC_4 VDD VDDI TSMC_7 VSS TSMC_9 TSMC_17 
+ S6ALLSVTFW8U20_RF_RXDEC 
XIXDEC<0> TSMC_16 TSMC_1 TSMC_6 VDD VDDI TSMC_7 VSS TSMC_11 TSMC_17 
+ S6ALLSVTFW8U20_RF_RXDEC 
XI64<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI64<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<3> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<2> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<1> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI65<0> TSMC_13 TSMC_12 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RXDECX4_LR
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RXDECX4_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI TSMC_7 VSS TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
XIXDEC_LR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDD VDDI TSMC_7 VSS 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 
+ S6ALLSVTFW8U20_RF_RXDECX4 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_XDEC4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_XDEC4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 VDD VDDI TSMC_42 VSS 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 
XXwdec TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 VDD VDDI TSMC_42 VSS 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_69 TSMC_70 
+ S6ALLSVTFW8U20_RF_WXDECX4_LR 
XXrdec TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 VDD VDDI TSMC_42 VSS 
+ TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_67 TSMC_68 
+ S6ALLSVTFW8U20_RF_RXDECX4_LR 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TIELGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TIELGEN TSMC_1 TSMC_2 VDD VSS 
MM5 TSMC_1 TSMC_2 VDD VDD pch_svt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_3 TSMC_4 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_2 TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=3 m=2 
MM2 TSMC_3 TSMC_5 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_2 TSMC_6 VSS VSS nch_svt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_3 TSMC_5 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI0 VSS VSS TSMC_5 TSMC_4 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI1 VSS VSS TSMC_4 TSMC_6 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PUDELAY
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_PUDELAY TSMC_1 TSMC_2 TSMC_3 VDD VSS 
XI3 VSS VSS TSMC_4 TSMC_2 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=5 n_l=0.020u p_totalM=3 p_nfin=5 p_l=0.020u 
XI149 TSMC_1 TSMC_3 VSS VSS VDD VDD TSMC_4 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DEC2TO4
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_DEC2TO4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS 
XI26 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI27 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI28 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI33 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI34 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI37 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI31 VSS VSS TSMC_10 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI35 VSS VSS TSMC_11 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI39 VSS VSS TSMC_12 TSMC_5 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI29 VSS VSS TSMC_9 TSMC_8 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_YDEC3TO8L
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_YDEC3TO8L TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
XI32 TSMC_3 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI42 TSMC_6 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI38 TSMC_6 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI43 TSMC_3 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI39 TSMC_3 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_19 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI35 TSMC_6 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_3 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_6 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 VSS VSS TSMC_17 TSMC_23 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI82 VSS VSS TSMC_24 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI15 VSS VSS TSMC_25 TSMC_14 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI85 VSS VSS TSMC_26 TSMC_9 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI3 VSS VSS TSMC_22 TSMC_25 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI94 VSS VSS TSMC_18 TSMC_27 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI93 VSS VSS TSMC_16 TSMC_28 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI81 VSS VSS TSMC_29 TSMC_13 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI87 VSS VSS TSMC_27 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI92 VSS VSS TSMC_19 TSMC_26 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI90 VSS VSS TSMC_21 TSMC_30 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI83 VSS VSS TSMC_30 TSMC_11 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI84 VSS VSS TSMC_23 TSMC_10 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
XI89 VSS VSS TSMC_20 TSMC_24 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI88 VSS VSS TSMC_15 TSMC_29 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=2 p_nfin=3 p_l=0.020u 
XI86 VSS VSS TSMC_28 TSMC_8 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.020u p_totalM=4 p_nfin=8 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DECPDA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_DECPDA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS 
XI58 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI60 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI59 TSMC_1 TSMC_4 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_3 TSMC_4 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI61 VSS VSS TSMC_9 TSMC_13 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI64 VSS VSS TSMC_11 TSMC_14 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI66 VSS VSS TSMC_15 TSMC_5 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI62 VSS VSS TSMC_13 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI63 VSS VSS TSMC_14 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI65 VSS VSS TSMC_10 TSMC_15 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI35 VSS VSS TSMC_16 TSMC_8 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=8 n_l=0.020u p_totalM=6 p_nfin=8 p_l=0.020u 
XI42 VSS VSS TSMC_12 TSMC_16 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RPREDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RPREDEC TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI VSS TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 
XXpb TSMC_5 TSMC_6 TSMC_13 TSMC_14 TSMC_27 TSMC_28 TSMC_29 TSMC_30 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DEC2TO4 
XXpd TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DEC2TO4 
XXpc TSMC_3 TSMC_4 TSMC_11 TSMC_12 TSMC_31 TSMC_32 TSMC_33 TSMC_34 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DEC2TO4 
XXya TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 VDD VDDI VSS TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ S6ALLSVTFW8U20_RF_YDEC3TO8L 
XXpa TSMC_7 TSMC_8 TSMC_15 TSMC_16 TSMC_23 TSMC_24 TSMC_25 TSMC_26 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DECPDA 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RPRCHBUF
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RPRCHBUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_1 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI43 VSS VSS TSMC_3 TSMC_7 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=6 n_l=0.020u p_totalM=3 p_nfin=4 p_l=0.020u 
XI42 VSS VSS TSMC_1 TSMC_2 TSMC_6 VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI2 VSS VSS TSMC_7 TSMC_4 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=13 n_nfin=5 n_l=0.020u p_totalM=13 p_nfin=9 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RCLKGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RCLKGEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS 
XI53 TSMC_11 TSMC_2 VSS VSS VDDI VDD TSMC_12 
+ S6ALLSVTFW8U20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=8 p_l=0.016u 
XI25 TSMC_13 TSMC_2 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nor2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
XI73 VSS VSS TSMC_9 TSMC_15 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI5 VSS VSS TSMC_13 TSMC_16 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI6 VSS VSS TSMC_13 TSMC_3 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=9 n_nfin=5 n_l=0.016u p_totalM=9 p_nfin=5 p_l=0.016u 
XI40 VSS VSS TSMC_12 TSMC_17 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI2 VSS VSS TSMC_18 TSMC_19 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI29 VSS VSS TSMC_2 TSMC_20 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI19 VSS VSS TSMC_1 TSMC_2 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI79 VSS VSS TSMC_7 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=2 n_nfin=5 n_l=0.016u p_totalM=2 p_nfin=5 p_l=0.016u 
XI17 VSS VSS TSMC_15 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=2 n_nfin=8 n_l=0.016u p_totalM=2 p_nfin=8 p_l=0.016u 
MM1 TSMC_21 TSMC_22 VDD VDD pch_ulvt_mac l=0.016u nfin=8 m=3 
MM3 TSMC_13 TSMC_4 TSMC_21 VDD pch_ulvt_mac l=0.016u nfin=8 m=3 
MM9 TSMC_18 TSMC_8 TSMC_23 VDD pch_ulvt_mac l=0.016u nfin=6 m=1 
MM5 TSMC_23 TSMC_20 VDDI VDD pch_ulvt_mac l=0.016u nfin=6 m=1 
MM13 TSMC_24 TSMC_12 VDD VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM6 TSMC_18 TSMC_19 TSMC_25 VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM12 TSMC_13 TSMC_16 TSMC_24 VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM10 TSMC_25 TSMC_14 VDDI VDD pch_ulvt_mac l=0.016u nfin=2 m=1 
MM0 TSMC_16 TSMC_8 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=2 
MM8 TSMC_13 TSMC_12 VSS VSS nch_ulvt_mac l=0.016u nfin=5 m=6 
MM4 TSMC_26 TSMC_20 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM11 TSMC_18 TSMC_8 VSS VSS nch_ulvt_mac l=0.016u nfin=4 m=1 
MM2 TSMC_18 TSMC_14 VSS VSS nch_ulvt_mac l=0.016u nfin=4 m=1 
MM15 TSMC_27 TSMC_16 VSS VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM7 TSMC_18 TSMC_19 TSMC_26 VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
MM14 TSMC_13 TSMC_16 TSMC_27 VSS nch_ulvt_mac l=0.016u nfin=2 m=1 
XI71 TSMC_13 TSMC_28 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nand2_ulvt_mac_pcell n_totalM=2 n_nfin=3 n_l=0.016u p_totalM=2 
+ p_nfin=3 p_l=0.016u 
XI75 TSMC_5 TSMC_20 VSS VSS VDD VDD TSMC_28 
+ S6ALLSVTFW8U20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI56 TSMC_18 TSMC_5 VSS VSS VDD VDD TSMC_11 
+ S6ALLSVTFW8U20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI82 TSMC_29 TSMC_17 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW8U20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
XI8 TSMC_20 TSMC_10 VSS VSS VDDI VDD TSMC_29 
+ S6ALLSVTFW8U20_nand2_ulvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH_RA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_ILATCH_RA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_ulvt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_ulvt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_ulvt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW8U20_inv_ulvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_ulvt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_ulvt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_ulvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH_RA_Y
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_ILATCH_RA_Y TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI 
+ VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_lvt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_lvt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_lvt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW8U20_inv_lvt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_lvt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_lvt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ADRLAT_RA
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_ADRLAT_RA TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 VDD VDDI VSS 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 
XXxlat<7> TSMC_25 TSMC_1 TSMC_2 TSMC_3 TSMC_11 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXxlat<6> TSMC_26 TSMC_1 TSMC_2 TSMC_4 TSMC_12 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXxlat<5> TSMC_27 TSMC_1 TSMC_2 TSMC_5 TSMC_13 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXxlat<4> TSMC_28 TSMC_1 TSMC_2 TSMC_6 TSMC_14 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXxlat<3> TSMC_29 TSMC_1 TSMC_2 TSMC_7 TSMC_15 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXxlat<2> TSMC_30 TSMC_1 TSMC_2 TSMC_8 TSMC_16 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXxlat<1> TSMC_31 TSMC_1 TSMC_2 TSMC_9 TSMC_17 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXxlat<0> TSMC_32 TSMC_1 TSMC_2 TSMC_10 TSMC_18 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA 
XXylat<2> TSMC_33 TSMC_1 TSMC_2 TSMC_19 TSMC_22 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA_Y 
XXylat<1> TSMC_34 TSMC_1 TSMC_2 TSMC_20 TSMC_23 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA_Y 
XXylat<0> TSMC_35 TSMC_1 TSMC_2 TSMC_21 TSMC_24 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH_RA_Y 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RENLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RENLAT TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
XI15 VSS VSS TSMC_5 TSMC_3 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI0 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI5 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
MM4 TSMC_8 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_9 TSMC_5 TSMC_8 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_10 TSMC_6 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_9 TSMC_2 TSMC_10 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_9 TSMC_5 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_11 TSMC_6 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_9 TSMC_2 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_12 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI6 TSMC_4 TSMC_9 VSS VSS VDD VDD TSMC_5 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RTUNE
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RTUNE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDI VSS 
XXenlat TSMC_1 TSMC_10 TSMC_8 TSMC_9 VDD VDDI VSS 
+ S6ALLSVTFW8U20_RF_RENLAT 
XI12<2> VSS VSS TSMC_13 TSMC_5 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI12<1> VSS VSS TSMC_14 TSMC_6 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI12<0> VSS VSS TSMC_15 TSMC_7 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=5 p_l=0.020u 
XI13<2> VSS VSS TSMC_2 TSMC_13 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI13<1> VSS VSS TSMC_3 TSMC_14 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI13<0> VSS VSS TSMC_4 TSMC_15 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI7 VSS VSS TSMC_11 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=5 n_l=0.020u p_totalM=4 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RGCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RGCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 VDD VDDI VSS TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
XXpredecs TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
+ TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 VDD VDDI VSS TSMC_58 
+ TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ S6ALLSVTFW8U20_RF_RPREDEC 
XXrprchb TSMC_38 TSMC_82 TSMC_83 TSMC_43 TSMC_46 VDD VDDI VSS 
+ S6ALLSVTFW8U20_RF_RPRCHBUF 
XXclkgen TSMC_1 TSMC_84 TSMC_40 TSMC_44 TSMC_85 TSMC_8 TSMC_9 TSMC_38 TSMC_83 
+ TSMC_45 VDD VDDI VSS S6ALLSVTFW8U20_RF_RCLKGEN 
XXadrlat TSMC_8 TSMC_9 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 VDD VDDI VSS 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 S6ALLSVTFW8U20_RF_ADRLAT_RA 
XXrtune TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_85 
+ TSMC_82 TSMC_39 TSMC_41 TSMC_42 VDD VDDI VSS S6ALLSVTFW8U20_RF_RTUNE 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_DKCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_DKCTD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI VSS 
MM2 VDDI TSMC_5 VDDI VDD pch_svt_mac l=0.020u nfin=4 m=1 
MM1 VSS TSMC_5 VSS VSS nch_svt_mac l=0.020u nfin=4 m=1 
XI126 TSMC_4 TSMC_5 VSS VSS VDDI VDD TSMC_6 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=2 n_nfin=2 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI64 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_7 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI76 TSMC_8 TSMC_9 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 
+ p_nfin=4 p_l=0.020u 
XI66 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_11 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_12 TSMC_6 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI179 TSMC_14 TSMC_6 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI178 TSMC_16 TSMC_6 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_1 TSMC_18 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_2 TSMC_19 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI156 TSMC_6 TSMC_10 VSS VSS VDDI VDD TSMC_3 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=6 n_nfin=10 n_l=0.020u p_totalM=6 
+ p_nfin=5 p_l=0.020u 
XI89 VSS VSS TSMC_11 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_7 TSMC_8 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_15 TSMC_20 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_21 TSMC_19 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_17 TSMC_22 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_20 TSMC_18 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_22 TSMC_9 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_13 TSMC_21 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WCLKGEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WCLKGEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS TSMC_9 
MM11 TSMC_10 TSMC_11 TSMC_12 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM10 TSMC_12 TSMC_13 VDDI VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM13 TSMC_14 TSMC_15 VDD VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM2 TSMC_16 TSMC_17 VDDI VDD pch_svt_mac l=0.016u nfin=6 m=1 
MM3 TSMC_18 TSMC_3 TSMC_19 VDD pch_svt_mac l=0.016u nfin=8 m=3 
MM1 TSMC_19 TSMC_20 VDD VDD pch_svt_mac l=0.016u nfin=8 m=3 
MM0 TSMC_10 TSMC_7 TSMC_16 VDD pch_svt_mac l=0.016u nfin=6 m=1 
MM12 TSMC_18 TSMC_21 TSMC_14 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM15 TSMC_22 TSMC_21 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM7 TSMC_10 TSMC_11 TSMC_23 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM14 TSMC_18 TSMC_21 TSMC_22 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM4 TSMC_23 TSMC_17 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM9 TSMC_21 TSMC_7 VSS VSS nch_svt_mac l=0.016u nfin=2 m=2 
MM8 TSMC_18 TSMC_15 VSS VSS nch_svt_mac l=0.016u nfin=5 m=6 
MM5 TSMC_10 TSMC_7 VSS VSS nch_svt_mac l=0.016u nfin=4 m=1 
MM6 TSMC_10 TSMC_13 VSS VSS nch_svt_mac l=0.016u nfin=4 m=1 
XI61 VSS VSS TSMC_24 TSMC_9 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=5 n_l=0.016u p_totalM=6 p_nfin=5 p_l=0.016u 
XI48 VSS VSS TSMC_18 TSMC_6 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=8 n_l=0.016u p_totalM=3 p_nfin=9 p_l=0.016u 
XI45 VSS VSS TSMC_18 TSMC_25 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI28 VSS VSS TSMC_26 TSMC_24 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=8 n_l=0.016u p_totalM=1 p_nfin=8 p_l=0.016u 
XI17 VSS VSS TSMC_6 TSMC_5 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=8 n_l=0.016u p_totalM=1 p_nfin=8 p_l=0.016u 
XI44 VSS VSS TSMC_25 TSMC_27 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.016u p_totalM=2 p_nfin=4 p_l=0.016u 
XI5 VSS VSS TSMC_18 TSMC_21 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI29 VSS VSS TSMC_18 TSMC_26 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI6 VSS VSS TSMC_27 TSMC_2 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=6 n_nfin=5 n_l=0.016u p_totalM=6 p_nfin=5 p_l=0.016u 
XI26 VSS VSS TSMC_24 TSMC_9 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=8 n_l=0.016u p_totalM=4 p_nfin=8 p_l=0.016u 
XI2 VSS VSS TSMC_10 TSMC_11 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI1 VSS VSS TSMC_28 TSMC_17 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI0 VSS VSS TSMC_1 TSMC_28 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 p_nfin=4 p_l=0.016u 
XI40 VSS VSS TSMC_15 TSMC_29 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
XI8 TSMC_17 TSMC_8 VSS VSS VDDI VDD TSMC_30 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI37 TSMC_30 TSMC_29 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
XI52 TSMC_10 TSMC_4 VSS VSS VDD VDD TSMC_31 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=2 p_l=0.016u 
XI53 TSMC_31 TSMC_28 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=4 n_l=0.016u p_totalM=1 
+ p_nfin=8 p_l=0.016u 
XI50 TSMC_18 TSMC_28 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 
+ p_nfin=3 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_YDEC3TO8
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_YDEC3TO8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDD VDDI VSS TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
XI32 TSMC_3 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_15 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI35 TSMC_6 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_16 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI36 TSMC_3 TSMC_2 TSMC_4 VSS VSS VDDI VDD TSMC_17 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI38 TSMC_6 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_18 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI39 TSMC_3 TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_19 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI42 TSMC_6 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI43 TSMC_3 TSMC_2 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI55 TSMC_6 TSMC_5 TSMC_4 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI33 VSS VSS TSMC_15 TSMC_13 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI34 VSS VSS TSMC_16 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI37 VSS VSS TSMC_17 TSMC_11 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI40 VSS VSS TSMC_18 TSMC_10 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI41 VSS VSS TSMC_19 TSMC_9 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI44 VSS VSS TSMC_20 TSMC_8 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI29 VSS VSS TSMC_22 TSMC_14 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
XI45 VSS VSS TSMC_21 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=3 n_l=0.020u p_totalM=1 p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WPREDEC
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WPREDEC TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI VSS TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 
XXya TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 VDD VDDI VSS TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ S6ALLSVTFW8U20_RF_YDEC3TO8 
XXpb TSMC_5 TSMC_6 TSMC_13 TSMC_14 TSMC_27 TSMC_28 TSMC_29 TSMC_30 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DEC2TO4 
XXpd TSMC_1 TSMC_2 TSMC_9 TSMC_10 TSMC_35 TSMC_36 TSMC_37 TSMC_38 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DEC2TO4 
XXpc TSMC_3 TSMC_4 TSMC_11 TSMC_12 TSMC_31 TSMC_32 TSMC_33 TSMC_34 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DEC2TO4 
XXpa TSMC_7 TSMC_8 TSMC_15 TSMC_16 TSMC_23 TSMC_24 TSMC_25 TSMC_26 VDD VDDI 
+ VSS S6ALLSVTFW8U20_RF_DECPDA 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ENLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_ENLAT TSMC_1 TSMC_2 TSMC_3 VDD VDDI VSS 
XI0 VSS VSS TSMC_1 TSMC_4 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI6 VSS VSS TSMC_5 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI5 VSS VSS TSMC_4 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI4 VSS VSS TSMC_6 TSMC_3 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
MM5 TSMC_5 TSMC_6 TSMC_8 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_8 TSMC_7 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_5 TSMC_2 TSMC_9 VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_9 TSMC_4 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_5 TSMC_6 TSMC_10 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_10 TSMC_4 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_5 TSMC_2 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_11 TSMC_7 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WTUNE
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WTUNE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDI VSS TSMC_9 TSMC_10 TSMC_11 
XXenlat TSMC_1 TSMC_9 TSMC_8 VDD VDDI VSS S6ALLSVTFW8U20_RF_ENLAT 
XI15 VSS VSS TSMC_10 TSMC_11 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=3 n_nfin=7 n_l=0.020u p_totalM=3 p_nfin=7 p_l=0.020u 
XI9<2> VSS VSS TSMC_2 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI9<1> VSS VSS TSMC_3 TSMC_13 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI9<0> VSS VSS TSMC_4 TSMC_14 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI8<2> VSS VSS TSMC_12 TSMC_5 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 p_nfin=5 p_l=0.020u 
XI8<1> VSS VSS TSMC_13 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 p_nfin=5 p_l=0.020u 
XI8<0> VSS VSS TSMC_14 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WPRCHBUF
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WPRCHBUF TSMC_1 TSMC_2 VDD VDDI VSS TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
XI18 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_20 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=2 n_nfin=5 n_l=0.020u p_totalM=2 
+ p_nfin=7 p_l=0.020u 
XI17<7> TSMC_8 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<6> TSMC_9 TSMC_1 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<5> TSMC_10 TSMC_1 VSS VSS VDDI VDD TSMC_23 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<4> TSMC_11 TSMC_1 VSS VSS VDDI VDD TSMC_24 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<3> TSMC_4 TSMC_1 VSS VSS VDDI VDD TSMC_25 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<2> TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_26 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<1> TSMC_6 TSMC_1 VSS VSS VDDI VDD TSMC_27 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI17<0> TSMC_7 TSMC_1 VSS VSS VDDI VDD TSMC_28 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<7> TSMC_8 TSMC_1 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<6> TSMC_9 TSMC_1 VSS VSS VDDI VDD TSMC_22 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<5> TSMC_10 TSMC_1 VSS VSS VDDI VDD TSMC_23 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<4> TSMC_11 TSMC_1 VSS VSS VDDI VDD TSMC_24 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<3> TSMC_4 TSMC_1 VSS VSS VDDI VDD TSMC_25 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<2> TSMC_5 TSMC_1 VSS VSS VDDI VDD TSMC_26 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<1> TSMC_6 TSMC_1 VSS VSS VDDI VDD TSMC_27 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI9<0> TSMC_7 TSMC_1 VSS VSS VDDI VDD TSMC_28 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=5 n_l=0.020u p_totalM=1 
+ p_nfin=5 p_l=0.020u 
XI7<7> VSS VSS TSMC_21 TSMC_12 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<6> VSS VSS TSMC_22 TSMC_13 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<5> VSS VSS TSMC_23 TSMC_14 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<4> VSS VSS TSMC_24 TSMC_15 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<3> VSS VSS TSMC_25 TSMC_16 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<2> VSS VSS TSMC_26 TSMC_17 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<1> VSS VSS TSMC_27 TSMC_18 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI7<0> VSS VSS TSMC_28 TSMC_19 VDDI VDD 
+ S6ALLSVTFW8U20_inv_svt_mac_pcell n_totalM=4 n_nfin=9 n_l=0.020u p_totalM=4 
+ p_nfin=9 p_l=0.020u 
XI2 VSS VSS TSMC_20 TSMC_3 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=4 n_nfin=9 n_l=16.0n p_totalM=6 p_nfin=9 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    ILATCH
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_ILATCH TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDD VDDI VSS 
MM6 TSMC_6 TSMC_7 TSMC_8 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_8 TSMC_2 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_9 TSMC_3 VDDI VDD pch_svt_mac l=0.020u nfin=3 m=1 
MM1 TSMC_6 TSMC_1 TSMC_9 VDD pch_svt_mac l=0.020u nfin=3 m=1 
XI7 VSS VSS TSMC_6 TSMC_4 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
XI6 VSS VSS TSMC_6 TSMC_7 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI22 VSS VSS TSMC_7 TSMC_5 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=4 n_l=0.020u p_totalM=1 p_nfin=4 p_l=0.020u 
MM2 TSMC_6 TSMC_1 TSMC_10 VSS nch_svt_mac l=0.020u nfin=3 m=1 
MM3 TSMC_10 TSMC_2 VSS VSS nch_svt_mac l=0.020u nfin=3 m=1 
MM4 TSMC_11 TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MM5 TSMC_6 TSMC_7 TSMC_11 VSS nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_ADRLAT
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_ADRLAT TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 VDD VDDI VSS 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 
XXylat<2> TSMC_33 TSMC_1 TSMC_2 TSMC_19 TSMC_22 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXylat<1> TSMC_34 TSMC_1 TSMC_2 TSMC_20 TSMC_23 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXylat<0> TSMC_35 TSMC_1 TSMC_2 TSMC_21 TSMC_24 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<7> TSMC_25 TSMC_1 TSMC_2 TSMC_3 TSMC_11 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<6> TSMC_26 TSMC_1 TSMC_2 TSMC_4 TSMC_12 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<5> TSMC_27 TSMC_1 TSMC_2 TSMC_5 TSMC_13 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<4> TSMC_28 TSMC_1 TSMC_2 TSMC_6 TSMC_14 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<3> TSMC_29 TSMC_1 TSMC_2 TSMC_7 TSMC_15 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<2> TSMC_30 TSMC_1 TSMC_2 TSMC_8 TSMC_16 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<1> TSMC_31 TSMC_1 TSMC_2 TSMC_9 TSMC_17 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
XXxlat<0> TSMC_32 TSMC_1 TSMC_2 TSMC_10 TSMC_18 VDD VDDI VSS 
+ S6ALLSVTFW8U20_ILATCH 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WGCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WGCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 VDD VDDI VSS TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 
XXclkgen TSMC_1 TSMC_33 TSMC_38 TSMC_62 TSMC_8 TSMC_9 TSMC_26 TSMC_31 VDD VDDI 
+ VSS TSMC_36 S6ALLSVTFW8U20_RF_WCLKGEN 
XXpredecs TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 
+ TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_10 TSMC_11 
+ TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 VDD VDDI VSS TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ S6ALLSVTFW8U20_RF_WPREDEC 
XXwtune TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_62 VDD VDDI VSS 
+ TSMC_32 TSMC_34 TSMC_35 S6ALLSVTFW8U20_RF_WTUNE 
XXwprchb TSMC_9 TSMC_26 VDD VDDI VSS TSMC_37 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 S6ALLSVTFW8U20_RF_WPRCHBUF 
XXadrlat TSMC_8 TSMC_9 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 VDD VDDI VSS 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 S6ALLSVTFW8U20_RF_ADRLAT 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_GCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_GCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 VDD VDDI VSS TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 
+ TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 
XXtiel TSMC_87 TSMC_88 VDD VSS S6ALLSVTFW8U20_RF_TIELGEN 
XXpudelay TSMC_27 TSMC_30 TSMC_86 VDD VSS S6ALLSVTFW8U20_RF_PUDELAY 
XXrctrl TSMC_1 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_39 
+ TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_20 
+ TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_29 TSMC_35 TSMC_36 TSMC_37 
+ TSMC_38 TSMC_71 TSMC_73 TSMC_89 TSMC_90 VDD VDDI VSS TSMC_75 TSMC_76 
+ TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 
+ TSMC_85 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 S6ALLSVTFW8U20_RF_RGCTRL 
XXdkctd TSMC_8 TSMC_9 TSMC_3 TSMC_13 TSMC_7 VDD VDDI VSS 
+ S6ALLSVTFW8U20_RF_DKCTD 
XXwctrl TSMC_2 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_29 TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_89 VDD VDDI VSS 
+ TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 
+ TSMC_124 TSMC_125 TSMC_126 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 
+ S6ALLSVTFW8U20_RF_WGCTRL 
MM1_header VDDI TSMC_28 VDD VDD pch_svt_mac l=0.020u nfin=7 m=24 
XI13 VSS VSS TSMC_28 TSMC_139 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=4 n_l=0.020u p_totalM=2 p_nfin=4 p_l=0.020u 
XI29 VSS VSS TSMC_88 TSMC_140 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=6 n_l=0.020u p_totalM=1 p_nfin=6 p_l=0.020u 
XI3 VSS VSS TSMC_140 TSMC_141 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=2 n_nfin=6 n_l=0.020u p_totalM=2 p_nfin=6 p_l=0.020u 
XI12 VSS VSS TSMC_139 TSMC_29 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=8 n_nfin=5 n_l=0.020u p_totalM=8 p_nfin=5 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RCTD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RCTD TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI VSS 
XI79 TSMC_5 TSMC_6 VSS VSS VDDI VDD TSMC_7 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI90 TSMC_2 TSMC_8 VSS VSS VDDI VDD TSMC_9 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI78 TSMC_9 TSMC_6 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI76 TSMC_11 TSMC_10 VSS VSS VDDI VDD TSMC_4 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI86 TSMC_12 TSMC_6 VSS VSS VDDI VDD TSMC_13 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI66 TSMC_2 TSMC_3 VSS VSS VDDI VDD TSMC_14 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI91 TSMC_3 TSMC_15 VSS VSS VDDI VDD TSMC_5 
+ S6ALLSVTFW8U20_nand2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
XI149 VSS VSS TSMC_13 TSMC_16 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI147 VSS VSS TSMC_11 TSMC_17 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI89 VSS VSS TSMC_14 TSMC_12 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI152 VSS VSS TSMC_7 TSMC_18 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI154 VSS VSS TSMC_19 TSMC_20 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI153 VSS VSS TSMC_18 TSMC_8 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI65 VSS VSS TSMC_21 TSMC_11 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI155 VSS VSS TSMC_20 TSMC_15 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI145 VSS VSS TSMC_1 TSMC_6 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI146 VSS VSS TSMC_11 TSMC_22 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI144 VSS VSS TSMC_23 TSMC_24 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI150 VSS VSS TSMC_13 TSMC_25 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI10 VSS VSS TSMC_16 TSMC_23 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI143 VSS VSS TSMC_24 TSMC_19 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI64 TSMC_3 TSMC_2 VSS VSS VDDI VDD TSMC_21 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_RDTRKEN
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_RDTRKEN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDI VSS 
MM24 TSMC_11 TSMC_10 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM17 TSMC_4 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=4 m=4 
MM16 TSMC_4 TSMC_10 TSMC_12 VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM15 TSMC_12 TSMC_6 VSS VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM13 TSMC_3 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=3 m=2 
MM8 TSMC_2 TSMC_10 TSMC_13 VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM2 TSMC_1 TSMC_14 TSMC_15 VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM4 TSMC_15 TSMC_9 VSS VSS nch_svt_mac l=0.016u nfin=2 m=1 
MM9 TSMC_16 TSMC_5 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM7 TSMC_13 TSMC_1 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM10 TSMC_3 TSMC_10 TSMC_16 VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM23 TSMC_2 TSMC_11 VSS VSS nch_svt_mac l=0.016u nfin=3 m=1 
MM3 VDDI TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM30 TSMC_10 TSMC_11 VDD VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM27 TSMC_2 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM20 TSMC_17 TSMC_6 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM19 TSMC_4 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=6 
MM18 TSMC_4 TSMC_11 TSMC_17 VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM14 TSMC_3 TSMC_10 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=2 
MM26 TSMC_3 TSMC_11 TSMC_18 VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM5 TSMC_19 TSMC_14 VDDI VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM0 TSMC_1 TSMC_14 TSMC_19 VDD pch_svt_mac l=0.016u nfin=2 m=1 
MM29 TSMC_2 TSMC_11 TSMC_20 VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM28 TSMC_20 TSMC_1 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM25 TSMC_18 TSMC_5 VDDI VDD pch_svt_mac l=0.016u nfin=4 m=1 
MM1 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.016u nfin=5 m=2 
XI33 TSMC_7 TSMC_2 TSMC_9 VSS VSS VDDI VDD TSMC_8 
+ S6ALLSVTFW8U20_nand3_svt_mac_pcell n_totalM=2 n_nfin=6 n_l=0.016u p_totalM=2 
+ p_nfin=3 p_l=0.016u 
XI1 VSS VSS TSMC_1 TSMC_14 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.016u p_totalM=1 p_nfin=2 p_l=0.016u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKGIORD
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TRKGIORD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 VDD VDDI VSS TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
XXrctd TSMC_4 TSMC_8 TSMC_9 TSMC_34 VDD VDDI VSS S6ALLSVTFW8U20_RF_RCTD 
XI23 VSS VSS TSMC_35 TSMC_36 VDDI VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI33 VSS VSS TSMC_18 TSMC_35 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XXrdtrken TSMC_4 TSMC_1 TSMC_2 TSMC_3 TSMC_5 TSMC_6 TSMC_34 TSMC_19 TSMC_36 
+ TSMC_20 TSMC_21 VDD VDDI VSS S6ALLSVTFW8U20_RF_RDTRKEN 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    16FF_2P_D130_v0d2_x1_for_BL_trk
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk TSMC_1 TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 VDD VSS TSMC_6 TSMC_7 TSMC_8 
MNpg_rp TSMC_3 TSMC_5 TSMC_9 VSS nchpg_8trpsr_mac l=20n nfin=2 m=1 
MNpd_rp TSMC_9 TSMC_1 VSS VSS nchpd_8trpsr_mac l=20n nfin=2 m=1 
MNpg_R TSMC_6 TSMC_8 TSMC_10 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MNpd_R TSMC_10 TSMC_11 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpd_L TSMC_11 TSMC_1 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpg_L TSMC_7 VSS TSMC_11 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MPpu_R TSMC_12 TSMC_11 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
MPpu_L TSMC_11 TSMC_1 TSMC_2 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    16FF_2P_D130_v0d2_x1_for_BL_trk_x2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 TSMC_1 TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 VDD VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 
XI1 TSMC_1 TSMC_3 TSMC_4 TSMC_5 TSMC_7 VDD VSS TSMC_10 TSMC_11 TSMC_12 
+ S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk 
XI0 TSMC_1 TSMC_2 TSMC_4 TSMC_6 TSMC_8 VDD VSS TSMC_9 TSMC_11 TSMC_13 
+ S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RBL_TRK_4X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_D130_ARRAY_RBL_TRK_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 VDD VDDAI 
+ VSS TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 
XI4 VDDAI TSMC_22 TSMC_5 TSMC_6 TSMC_8 TSMC_9 TSMC_12 TSMC_13 VDD VSS 
+ TSMC_23 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
+ S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
XI5 VDDAI TSMC_4 TSMC_22 TSMC_6 TSMC_10 TSMC_11 VSS VSS VDD VSS TSMC_15 
+ TSMC_23 TSMC_17 TSMC_20 TSMC_21 
+ S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_WL_TRACK
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_WL_TRACK TSMC_1 VSS TSMC_2 TSMC_3 
MMRWL VSS TSMC_1 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MMWWL1 VSS TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
MMWWL0q VSS TSMC_3 VSS VSS nch_svt_mac l=0.020u nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RWL_TRK_X2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ VDD VDDAI VSS TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
XI4 TSMC_5 VSS TSMC_5 TSMC_12 S6ALLSVTFW8U20_RF_WL_TRACK 
XI5 TSMC_5 VSS TSMC_5 TSMC_12 S6ALLSVTFW8U20_RF_WL_TRACK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PIN_GCTRL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_PIN_GCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 VSS TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 
XD40 VSS TSMC_77 ndio_mac nfin=2 l=200.0n m=1 
XD39 VSS TSMC_49 ndio_mac nfin=2 l=200.0n m=1 
XD34 VSS TSMC_88 ndio_mac nfin=2 l=200.0n m=1 
XD41 VSS TSMC_78 ndio_mac nfin=2 l=200.0n m=1 
XD5<10> VSS TSMC_12 ndio_mac nfin=2 l=200.0n m=1 
XD5<9> VSS TSMC_13 ndio_mac nfin=2 l=200.0n m=1 
XD5<8> VSS TSMC_14 ndio_mac nfin=2 l=200.0n m=1 
XD5<7> VSS TSMC_15 ndio_mac nfin=2 l=200.0n m=1 
XD5<6> VSS TSMC_16 ndio_mac nfin=2 l=200.0n m=1 
XD5<5> VSS TSMC_17 ndio_mac nfin=2 l=200.0n m=1 
XD5<4> VSS TSMC_18 ndio_mac nfin=2 l=200.0n m=1 
XD5<3> VSS TSMC_19 ndio_mac nfin=2 l=200.0n m=1 
XD5<2> VSS TSMC_20 ndio_mac nfin=2 l=200.0n m=1 
XD5<1> VSS TSMC_21 ndio_mac nfin=2 l=200.0n m=1 
XD5<0> VSS TSMC_22 ndio_mac nfin=2 l=200.0n m=1 
XD8 VSS TSMC_81 ndio_mac nfin=2 l=200.0n m=1 
XD4<10> VSS TSMC_34 ndio_mac nfin=2 l=200.0n m=1 
XD4<9> VSS TSMC_35 ndio_mac nfin=2 l=200.0n m=1 
XD4<8> VSS TSMC_36 ndio_mac nfin=2 l=200.0n m=1 
XD4<7> VSS TSMC_37 ndio_mac nfin=2 l=200.0n m=1 
XD4<6> VSS TSMC_38 ndio_mac nfin=2 l=200.0n m=1 
XD4<5> VSS TSMC_39 ndio_mac nfin=2 l=200.0n m=1 
XD4<4> VSS TSMC_40 ndio_mac nfin=2 l=200.0n m=1 
XD4<3> VSS TSMC_41 ndio_mac nfin=2 l=200.0n m=1 
XD4<2> VSS TSMC_42 ndio_mac nfin=2 l=200.0n m=1 
XD4<1> VSS TSMC_43 ndio_mac nfin=2 l=200.0n m=1 
XD4<0> VSS TSMC_44 ndio_mac nfin=2 l=200.0n m=1 
XD25 VSS TSMC_48 ndio_mac nfin=2 l=200.0n m=1 
XD31<2> VSS TSMC_67 ndio_mac nfin=2 l=200.0n m=1 
XD31<1> VSS TSMC_68 ndio_mac nfin=2 l=200.0n m=1 
XD31<0> VSS TSMC_69 ndio_mac nfin=2 l=200.0n m=1 
XD21 VSS TSMC_92 ndio_mac nfin=2 l=200.0n m=1 
XD35<1> VSS TSMC_51 ndio_mac nfin=2 l=200.0n m=1 
XD35<0> VSS TSMC_52 ndio_mac nfin=2 l=200.0n m=1 
XDdummy<0> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<1> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<2> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<3> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<4> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XDdummy<5> VSS VSS ndio_mac nfin=2 l=200.0n m=1 
XD30<2> VSS TSMC_64 ndio_mac nfin=2 l=200.0n m=1 
XD30<1> VSS TSMC_65 ndio_mac nfin=2 l=200.0n m=1 
XD30<0> VSS TSMC_66 ndio_mac nfin=2 l=200.0n m=1 
XD28 VSS TSMC_47 ndio_mac nfin=2 l=200.0n m=1 
XD7 VSS TSMC_76 ndio_mac nfin=2 l=200.0n m=1 
XD2<10> VSS TSMC_23 ndio_mac nfin=2 l=200.0n m=1 
XD2<9> VSS TSMC_24 ndio_mac nfin=2 l=200.0n m=1 
XD2<8> VSS TSMC_25 ndio_mac nfin=2 l=200.0n m=1 
XD2<7> VSS TSMC_26 ndio_mac nfin=2 l=200.0n m=1 
XD2<6> VSS TSMC_27 ndio_mac nfin=2 l=200.0n m=1 
XD2<5> VSS TSMC_28 ndio_mac nfin=2 l=200.0n m=1 
XD2<4> VSS TSMC_29 ndio_mac nfin=2 l=200.0n m=1 
XD2<3> VSS TSMC_30 ndio_mac nfin=2 l=200.0n m=1 
XD2<2> VSS TSMC_31 ndio_mac nfin=2 l=200.0n m=1 
XD2<1> VSS TSMC_32 ndio_mac nfin=2 l=200.0n m=1 
XD2<0> VSS TSMC_33 ndio_mac nfin=2 l=200.0n m=1 
XD3<10> VSS TSMC_1 ndio_mac nfin=2 l=200.0n m=1 
XD3<9> VSS TSMC_2 ndio_mac nfin=2 l=200.0n m=1 
XD3<8> VSS TSMC_3 ndio_mac nfin=2 l=200.0n m=1 
XD3<7> VSS TSMC_4 ndio_mac nfin=2 l=200.0n m=1 
XD3<6> VSS TSMC_5 ndio_mac nfin=2 l=200.0n m=1 
XD3<5> VSS TSMC_6 ndio_mac nfin=2 l=200.0n m=1 
XD3<4> VSS TSMC_7 ndio_mac nfin=2 l=200.0n m=1 
XD3<3> VSS TSMC_8 ndio_mac nfin=2 l=200.0n m=1 
XD3<2> VSS TSMC_9 ndio_mac nfin=2 l=200.0n m=1 
XD3<1> VSS TSMC_10 ndio_mac nfin=2 l=200.0n m=1 
XD3<0> VSS TSMC_11 ndio_mac nfin=2 l=200.0n m=1 
XD0<1> VSS TSMC_71 ndio_mac nfin=2 l=200.0n m=1 
XD0<0> VSS TSMC_72 ndio_mac nfin=2 l=200.0n m=1 
XD24 VSS TSMC_46 ndio_mac nfin=2 l=200.0n m=1 
XD26 VSS TSMC_45 ndio_mac nfin=2 l=200.0n m=1 
XD6 VSS TSMC_50 ndio_mac nfin=2 l=200.0n m=1 
XD9 VSS TSMC_73 ndio_mac nfin=2 l=200.0n m=1 
XD20 VSS TSMC_91 ndio_mac nfin=2 l=200.0n m=1 
XD19 VSS TSMC_74 ndio_mac nfin=2 l=200.0n m=1 
XD38<8> VSS TSMC_53 ndio_mac nfin=2 l=200.0n m=1 
XD38<7> VSS TSMC_54 ndio_mac nfin=2 l=200.0n m=1 
XD38<6> VSS TSMC_55 ndio_mac nfin=2 l=200.0n m=1 
XD38<5> VSS TSMC_56 ndio_mac nfin=2 l=200.0n m=1 
XD38<4> VSS TSMC_57 ndio_mac nfin=2 l=200.0n m=1 
XD38<3> VSS TSMC_58 ndio_mac nfin=2 l=200.0n m=1 
XD38<2> VSS TSMC_59 ndio_mac nfin=2 l=200.0n m=1 
XD38<1> VSS TSMC_60 ndio_mac nfin=2 l=200.0n m=1 
XD38<0> VSS TSMC_61 ndio_mac nfin=2 l=200.0n m=1 
XD37 VSS TSMC_75 ndio_mac nfin=2 l=200.0n m=1 
XD42<1> VSS TSMC_79 ndio_mac nfin=2 l=200.0n m=1 
XD42<0> VSS TSMC_80 ndio_mac nfin=2 l=200.0n m=1 
XD1<1> VSS TSMC_89 ndio_mac nfin=2 l=200.0n m=1 
XD1<0> VSS TSMC_90 ndio_mac nfin=2 l=200.0n m=1 
XD29 VSS TSMC_87 ndio_mac nfin=2 l=200.0n m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    N16_2PRF_BITCELL
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_N16_2PRF_BITCELL TSMC_1 TSMC_2 TSMC_3 VDD VSS TSMC_4 
+ TSMC_5 TSMC_6 
MNpg_rp TSMC_2 TSMC_3 TSMC_7 VSS nchpg_8trpsr_mac l=20n nfin=2 m=1 
MNpd_rp TSMC_7 TSMC_8 VSS VSS nchpd_8trpsr_mac l=20n nfin=2 m=1 
MNpd_L TSMC_9 TSMC_8 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpd_R TSMC_8 TSMC_9 VSS VSS nchpd_8tsr_mac l=20n nfin=2 m=1 
MNpg_R TSMC_5 TSMC_6 TSMC_8 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MNpg_L TSMC_4 TSMC_6 TSMC_9 VSS nchpg_8tsr_mac l=20n nfin=2 m=1 
MPpu_L TSMC_9 TSMC_8 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
MPpu_R TSMC_8 TSMC_9 TSMC_1 VDD pchpu_8tsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_4X2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_D130_ARRAY_4X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 VDD VDDAI VSS TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 
XI7 VDDAI TSMC_3 TSMC_7 VDD VSS TSMC_9 TSMC_11 TSMC_15 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
XI6 VDDAI TSMC_4 TSMC_8 VDD VSS TSMC_10 TSMC_12 TSMC_16 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
XI5 VDDAI TSMC_3 TSMC_8 VDD VSS TSMC_9 TSMC_11 TSMC_16 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
XI4 VDDAI TSMC_4 TSMC_7 VDD VSS TSMC_10 TSMC_12 TSMC_15 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
XI3 VDDAI TSMC_4 TSMC_6 VDD VSS TSMC_10 TSMC_12 TSMC_14 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
XI2 VDDAI TSMC_3 TSMC_6 VDD VSS TSMC_9 TSMC_11 TSMC_14 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
XI1 VDDAI TSMC_4 TSMC_5 VDD VSS TSMC_10 TSMC_12 TSMC_13 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
XI0 VDDAI TSMC_3 TSMC_5 VDD VSS TSMC_9 TSMC_11 TSMC_13 
+ S6ALLSVTFW8U20_N16_2PRF_BITCELL 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RBL_TRK_OFF_4X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_D130_ARRAY_RBL_TRK_OFF_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDD VDDAI VSS TSMC_12 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 
XI2 VDDAI TSMC_4 TSMC_20 TSMC_6 TSMC_10 TSMC_11 VSS VSS VDD VSS TSMC_12 
+ TSMC_21 TSMC_15 TSMC_18 TSMC_19 
+ S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
XI4 VDDAI TSMC_20 TSMC_5 TSMC_6 TSMC_8 TSMC_9 VSS VSS VDD VSS TSMC_21 
+ TSMC_13 TSMC_15 TSMC_16 TSMC_17 
+ S6ALLSVTFW8U20_16FF_2P_D130_v0d2_x1_for_BL_trk_x2 
.ENDS

************************************************************************
* Library Name: tsn16ff2prf_demo_array_d130
* Cell Name:    D130_ARRAY_RWL_TRK_X1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X1 TSMC_1 TSMC_2 TSMC_3 VDD VDDAI VSS 
+ TSMC_4 TSMC_5 TSMC_6 TSMC_7 
XI2 TSMC_3 VSS TSMC_3 TSMC_7 S6ALLSVTFW8U20_RF_WL_TRACK 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_PIN_GIO_MUX1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VSS 
XD3<1> VSS TSMC_3 ndio_mac nfin=2 l=200.0n m=1 
XD3<0> VSS TSMC_4 ndio_mac nfin=2 l=200.0n m=1 
XD2<1> VSS TSMC_1 ndio_mac nfin=2 l=200.0n m=1 
XD2<0> VSS TSMC_2 ndio_mac nfin=2 l=200.0n m=1 
XD0<1> VSS TSMC_5 ndio_mac nfin=2 l=200.0n m=1 
XD0<0> VSS TSMC_6 ndio_mac nfin=2 l=200.0n m=1 
XD1<1> VSS TSMC_7 ndio_mac nfin=2 l=200.0n m=1 
XD1<0> VSS TSMC_8 ndio_mac nfin=2 l=200.0n m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    LIO_PWR_TK_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_LIO_PWR_TK_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI 
+ TSMC_5 
MM_TKPKP3 TSMC_6 TSMC_3 TSMC_7 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP2 TSMC_7 TSMC_3 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP4 TSMC_5 TSMC_4 TSMC_6 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_TKPKP1 TSMC_6 TSMC_2 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKLIO_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TRKLIO_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDD VDDI VSS 
MM0 TSMC_3 TSMC_4 VSS VSS nch_lvt_mac l=0.020u nfin=7 m=2 
MM5 TSMC_11 TSMC_9 VSS VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM6 TSMC_1 TSMC_9 TSMC_11 VSS nch_lvt_mac l=0.020u nfin=2 m=1 
MM4 TSMC_9 TSMC_1 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM8 TSMC_12 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM2 TSMC_9 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=2 
MM11 VDD TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_9 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=2 
MM7 TSMC_14 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM13 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM14 TSMC_1 TSMC_9 VDDI VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_9 TSMC_1 TSMC_14 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI13 TSMC_5 TSMC_6 TSMC_7 TSMC_10 VDD VDDI TSMC_13 
+ S6ALLSVTFW8U20_LIO_PWR_TK_SVT_V1 
XXpwd0 TSMC_5 TSMC_6 TSMC_7 TSMC_10 VDD VDDI TSMC_13 
+ S6ALLSVTFW8U20_LIO_PWR_TK_SVT_V1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_TRKLIOX2_72_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_TRKLIOX2_72_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 VDD VDDAI VDDI VSS TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_23 TSMC_24 
XI35 VSS VSS TSMC_25 TSMC_26 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XI31 VSS VSS TSMC_27 TSMC_28 VDD VDD S6ALLSVTFW8U20_inv_svt_mac_pcell 
+ n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 p_nfin=2 p_l=0.020u 
XXtrklio TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_9 TSMC_10 TSMC_11 TSMC_26 TSMC_15 
+ TSMC_18 VDD VDDI VSS S6ALLSVTFW8U20_RF_TRKLIO_SVT_V1 
XI32 TSMC_14 TSMC_1 VSS VSS VDD VDD TSMC_27 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
XI38 TSMC_28 TSMC_16 VSS VSS VDD VDD TSMC_25 
+ S6ALLSVTFW8U20_nor2_svt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=3 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    LIO_PWR_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_LIO_PWR_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDD VDDI 
+ TSMC_5 
MM_PKP3 TSMC_5 TSMC_2 TSMC_6 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_PKP2 TSMC_6 TSMC_2 TSMC_7 VDD pch_svt_mac l=72.0n nfin=2 m=1 
MM_PKP1 TSMC_7 TSMC_2 VDD VDD pch_svt_mac l=72.0n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LIO_SVT_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_LIO_SVT_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 VDD VDDI VSS 
MM4 TSMC_1 TSMC_10 TSMC_11 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM8 TSMC_11 TSMC_8 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM3 TSMC_1 TSMC_7 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM0 TSMC_2 TSMC_8 VDD VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM1 TSMC_2 TSMC_10 TSMC_13 VDD pch_svt_mac l=0.020u nfin=2 m=1 
MM7 TSMC_13 TSMC_7 TSMC_12 VDD pch_svt_mac l=0.020u nfin=2 m=1 
XI0 TSMC_4 TSMC_5 TSMC_6 TSMC_9 VDD VDD TSMC_12 
+ S6ALLSVTFW8U20_LIO_PWR_SVT_V1 
MM2 TSMC_3 TSMC_10 VSS VSS nch_lvt_mac l=0.020u nfin=7 m=2 
XI17 TSMC_1 TSMC_2 VSS VSS VDDI VDD TSMC_10 
+ S6ALLSVTFW8U20_nand2_lvt_mac_pcell n_totalM=1 n_nfin=2 n_l=0.020u p_totalM=1 
+ p_nfin=2 p_l=0.020u 
.ENDS

************************************************************************
* Library Name: TS16FF2PRF
* Cell Name:    RF_LIOX2_72_V1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_RF_LIOX2_72_V1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDD VDDAI VDDI VSS TSMC_13 
+ TSMC_14 TSMC_15 TSMC_16 
XXlio0 TSMC_9 TSMC_11 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_12 
+ VDD VDDI VSS S6ALLSVTFW8U20_RF_LIO_SVT_V1 
XXlio1 TSMC_8 TSMC_10 TSMC_1 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_12 
+ VDD VDDI VSS S6ALLSVTFW8U20_RF_LIO_SVT_V1 
.ENDS

.SUBCKT ndio_mac PLUS MINUS 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_inv_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_ulvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_inv_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand3_ulvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nand3_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_lvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nor2_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nor2_ulvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nor2_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_lvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nand2_lvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    nand2_ulvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S6ALLSVTFW8U20_nand2_ulvt_mac_pcell TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS





**** End of leaf cells

.SUBCKT S6ALLSVTFW8U20_PIN_ROW TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 
+ TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 
+ TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 
+ TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 
+ TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 
+ TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 
+ TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 
+ TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 
+ TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 
+ TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 
+ TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 
+ TSMC_235 VSS TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_250 
XPINIO0 TSMC_95 TSMC_96 TSMC_209 TSMC_210 TSMC_31 TSMC_32 TSMC_177 TSMC_178 
+ TSMC_63 TSMC_64 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO1 TSMC_93 TSMC_94 TSMC_207 TSMC_208 TSMC_29 TSMC_30 TSMC_175 TSMC_176 
+ TSMC_61 TSMC_62 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO2 TSMC_91 TSMC_92 TSMC_205 TSMC_206 TSMC_27 TSMC_28 TSMC_173 TSMC_174 
+ TSMC_59 TSMC_60 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO3 TSMC_89 TSMC_90 TSMC_203 TSMC_204 TSMC_25 TSMC_26 TSMC_171 TSMC_172 
+ TSMC_57 TSMC_58 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO4 TSMC_87 TSMC_88 TSMC_201 TSMC_202 TSMC_23 TSMC_24 TSMC_169 TSMC_170 
+ TSMC_55 TSMC_56 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO5 TSMC_85 TSMC_86 TSMC_199 TSMC_200 TSMC_21 TSMC_22 TSMC_167 TSMC_168 
+ TSMC_53 TSMC_54 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO6 TSMC_83 TSMC_84 TSMC_197 TSMC_198 TSMC_19 TSMC_20 TSMC_165 TSMC_166 
+ TSMC_51 TSMC_52 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO7 TSMC_81 TSMC_82 TSMC_195 TSMC_196 TSMC_17 TSMC_18 TSMC_163 TSMC_164 
+ TSMC_49 TSMC_50 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO8 TSMC_79 TSMC_80 TSMC_193 TSMC_194 TSMC_15 TSMC_16 TSMC_161 TSMC_162 
+ TSMC_47 TSMC_48 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO9 TSMC_77 TSMC_78 TSMC_191 TSMC_192 TSMC_13 TSMC_14 TSMC_159 TSMC_160 
+ TSMC_45 TSMC_46 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO10 TSMC_75 TSMC_76 TSMC_189 TSMC_190 TSMC_11 TSMC_12 TSMC_157 TSMC_158 
+ TSMC_43 TSMC_44 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO11 TSMC_73 TSMC_74 TSMC_187 TSMC_188 TSMC_9 TSMC_10 TSMC_155 TSMC_156 
+ TSMC_41 TSMC_42 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO12 TSMC_71 TSMC_72 TSMC_185 TSMC_186 TSMC_7 TSMC_8 TSMC_153 TSMC_154 
+ TSMC_39 TSMC_40 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO13 TSMC_69 TSMC_70 TSMC_183 TSMC_184 TSMC_5 TSMC_6 TSMC_151 TSMC_152 
+ TSMC_37 TSMC_38 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO14 TSMC_67 TSMC_68 TSMC_181 TSMC_182 TSMC_3 TSMC_4 TSMC_149 TSMC_150 
+ TSMC_35 TSMC_36 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINIO15 TSMC_65 TSMC_66 TSMC_179 TSMC_180 TSMC_1 TSMC_2 TSMC_147 TSMC_148 
+ TSMC_33 TSMC_34 TSMC_251 TSMC_252 VSS 
+ S6ALLSVTFW8U20_RF_PIN_GIO_MUX1 
XPINCTRL TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 
+ TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_97 TSMC_98 TSMC_99 TSMC_100 
+ TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_211 TSMC_212 TSMC_213 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_136 
+ TSMC_235 TSMC_108 TSMC_121 TSMC_243 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 
+ TSMC_144 TSMC_145 TSMC_253 TSMC_254 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_236 TSMC_129 TSMC_130 TSMC_109 
+ TSMC_233 TSMC_146 TSMC_135 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_134 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_133 VSS TSMC_237 
+ TSMC_131 TSMC_132 TSMC_122 TSMC_234 S6ALLSVTFW8U20_RF_PIN_GCTRL 
.ENDS

.SUBCKT S6ALLSVTFW8U20_GCTRL_GIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 VDDI VDDM VSS TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 
+ TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 
+ TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 
+ TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 
+ TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 
+ TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 TSMC_344 
+ TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 
+ TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 
+ TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 TSMC_376 
+ TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 
+ TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 
+ TSMC_393 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 
+ TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 TSMC_408 
+ TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 
+ TSMC_417 TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 
+ TSMC_425 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 
+ TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 TSMC_440 
+ TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 
+ TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 
+ TSMC_457 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 
+ TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 TSMC_472 
+ TSMC_473 TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 
+ TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 
XGIO_MUX0 TSMC_33 TSMC_34 TSMC_65 TSMC_66 TSMC_97 TSMC_98 TSMC_488 TSMC_145 
+ TSMC_146 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_357 TSMC_358 TSMC_422 
+ TSMC_390 TSMC_218 TSMC_219 TSMC_250 TSMC_251 TSMC_285 TSMC_286 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX1 TSMC_31 TSMC_32 TSMC_63 TSMC_64 TSMC_95 TSMC_96 TSMC_488 TSMC_143 
+ TSMC_144 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_355 TSMC_356 TSMC_421 
+ TSMC_389 TSMC_216 TSMC_217 TSMC_248 TSMC_249 TSMC_283 TSMC_284 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX2 TSMC_29 TSMC_30 TSMC_61 TSMC_62 TSMC_93 TSMC_94 TSMC_488 TSMC_141 
+ TSMC_142 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_353 TSMC_354 TSMC_420 
+ TSMC_388 TSMC_214 TSMC_215 TSMC_246 TSMC_247 TSMC_281 TSMC_282 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX3 TSMC_27 TSMC_28 TSMC_59 TSMC_60 TSMC_91 TSMC_92 TSMC_488 TSMC_139 
+ TSMC_140 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_351 TSMC_352 TSMC_419 
+ TSMC_387 TSMC_212 TSMC_213 TSMC_244 TSMC_245 TSMC_279 TSMC_280 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX4 TSMC_25 TSMC_26 TSMC_57 TSMC_58 TSMC_89 TSMC_90 TSMC_488 TSMC_137 
+ TSMC_138 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_349 TSMC_350 TSMC_418 
+ TSMC_386 TSMC_210 TSMC_211 TSMC_242 TSMC_243 TSMC_277 TSMC_278 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX5 TSMC_23 TSMC_24 TSMC_55 TSMC_56 TSMC_87 TSMC_88 TSMC_488 
+ TSMC_135 TSMC_136 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_347 TSMC_348 TSMC_417 
+ TSMC_385 TSMC_208 TSMC_209 TSMC_240 TSMC_241 TSMC_275 TSMC_276 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX6 TSMC_21 TSMC_22 TSMC_53 TSMC_54 TSMC_85 TSMC_86 TSMC_488 
+ TSMC_133 TSMC_134 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_345 TSMC_346 TSMC_416 
+ TSMC_384 TSMC_206 TSMC_207 TSMC_238 TSMC_239 TSMC_273 TSMC_274 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX7 TSMC_19 TSMC_20 TSMC_51 TSMC_52 TSMC_83 TSMC_84 TSMC_488 
+ TSMC_131 TSMC_132 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_343 TSMC_344 TSMC_415 
+ TSMC_383 TSMC_204 TSMC_205 TSMC_236 TSMC_237 TSMC_271 TSMC_272 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX8 TSMC_17 TSMC_18 TSMC_49 TSMC_50 TSMC_81 TSMC_82 TSMC_488 
+ TSMC_129 TSMC_130 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_341 TSMC_342 TSMC_414 
+ TSMC_382 TSMC_202 TSMC_203 TSMC_234 TSMC_235 TSMC_269 TSMC_270 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX9 TSMC_15 TSMC_16 TSMC_47 TSMC_48 TSMC_79 TSMC_80 TSMC_488 
+ TSMC_127 TSMC_128 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_339 TSMC_340 TSMC_413 
+ TSMC_381 TSMC_200 TSMC_201 TSMC_232 TSMC_233 TSMC_267 TSMC_268 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX10 TSMC_13 TSMC_14 TSMC_45 TSMC_46 TSMC_77 TSMC_78 TSMC_488 
+ TSMC_125 TSMC_126 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_337 TSMC_338 TSMC_412 
+ TSMC_380 TSMC_198 TSMC_199 TSMC_230 TSMC_231 TSMC_265 TSMC_266 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX11 TSMC_11 TSMC_12 TSMC_43 TSMC_44 TSMC_75 TSMC_76 TSMC_488 
+ TSMC_123 TSMC_124 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_335 TSMC_336 TSMC_411 
+ TSMC_379 TSMC_196 TSMC_197 TSMC_228 TSMC_229 TSMC_263 TSMC_264 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX12 TSMC_9 TSMC_10 TSMC_41 TSMC_42 TSMC_73 TSMC_74 TSMC_488 
+ TSMC_121 TSMC_122 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_333 TSMC_334 TSMC_410 
+ TSMC_378 TSMC_194 TSMC_195 TSMC_226 TSMC_227 TSMC_261 TSMC_262 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX13 TSMC_7 TSMC_8 TSMC_39 TSMC_40 TSMC_71 TSMC_72 TSMC_488 
+ TSMC_119 TSMC_120 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_331 TSMC_332 TSMC_409 
+ TSMC_377 TSMC_192 TSMC_193 TSMC_224 TSMC_225 TSMC_259 TSMC_260 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX14 TSMC_5 TSMC_6 TSMC_37 TSMC_38 TSMC_69 TSMC_70 TSMC_488 
+ TSMC_117 TSMC_118 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_329 TSMC_330 TSMC_408 
+ TSMC_376 TSMC_190 TSMC_191 TSMC_222 TSMC_223 TSMC_257 TSMC_258 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_GIOM1X2 
XGIO_MUX15 TSMC_3 TSMC_4 TSMC_35 TSMC_36 TSMC_67 TSMC_68 TSMC_488 
+ TSMC_115 TSMC_116 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_327 TSMC_328 TSMC_407 
+ TSMC_375 TSMC_188 TSMC_189 TSMC_220 TSMC_221 TSMC_255 TSMC_256 
+ TSMC_490 TSMC_322 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_491 
+ TSMC_492 S6ALLSVTFW8U20_RF_GIOM1X2 
XTRKGIOL TSMC_488 TSMC_495 TSMC_496 TSMC_497 TSMC_498 TSMC_499 TSMC_500 
+ TSMC_501 TSMC_502 TSMC_489 TSMC_184 VDDM VDDI VSS TSMC_503 TSMC_504 
+ TSMC_112 TSMC_252 TSMC_253 TSMC_113 TSMC_490 TSMC_322 TSMC_505 
+ TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_491 TSMC_492 TSMC_493 
+ TSMC_494 S6ALLSVTFW8U20_RF_TRKGIOWR 
XTRKGIOR TSMC_510 TSMC_511 TSMC_512 TSMC_99 TSMC_185 TSMC_185 TSMC_488 TSMC_147 
+ TSMC_148 TSMC_495 TSMC_496 TSMC_497 TSMC_498 TSMC_499 TSMC_500 
+ TSMC_501 TSMC_502 TSMC_489 TSMC_513 TSMC_185 TSMC_184 VDDM VDDI VSS 
+ TSMC_319 TSMC_514 TSMC_490 TSMC_322 TSMC_506 TSMC_507 TSMC_508 
+ TSMC_509 TSMC_491 TSMC_492 TSMC_493 TSMC_494 
+ S6ALLSVTFW8U20_RF_TRKGIORD 
XGCTRL TSMC_1 TSMC_2 TSMC_324 TSMC_515 TSMC_325 TSMC_326 TSMC_323 TSMC_100 
+ TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 
+ TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_184 TSMC_184 TSMC_184 
+ TSMC_185 TSMC_185 TSMC_185 TSMC_516 TSMC_320 TSMC_114 TSMC_488 TSMC_321 
+ TSMC_185 TSMC_185 TSMC_185 TSMC_185 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_517 TSMC_518 TSMC_519 TSMC_520 
+ TSMC_521 TSMC_522 TSMC_495 TSMC_496 TSMC_497 TSMC_498 TSMC_499 TSMC_500 
+ TSMC_501 TSMC_502 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 
+ TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_489 TSMC_171 TSMC_513 
+ TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 
+ TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_487 TSMC_185 TSMC_184 
+ TSMC_186 TSMC_187 VDDM VDDI VSS TSMC_254 TSMC_287 TSMC_288 TSMC_289 
+ TSMC_490 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 
+ TSMC_296 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_322 TSMC_505 TSMC_308 
+ TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 TSMC_314 TSMC_315 
+ TSMC_316 TSMC_317 TSMC_318 TSMC_506 TSMC_507 TSMC_508 TSMC_509 
+ TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_523 TSMC_524 TSMC_525 
+ TSMC_526 S6ALLSVTFW8U20_RF_GCTRL 
.ENDS

.SUBCKT S6ALLSVTFW8U20_ROW_TRACKING TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 VDDM 
+ VDDAI VDDI VSS TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 
XTRKROW0 TSMC_95 TSMC_96 TSMC_104 TSMC_105 TSMC_101 VDDM VDDAI VSS TSMC_31 
+ TSMC_32 TSMC_63 TSMC_64 TSMC_106 TSMC_107 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW1 TSMC_93 TSMC_94 TSMC_108 TSMC_109 TSMC_101 VDDM VDDAI VSS TSMC_29 
+ TSMC_30 TSMC_61 TSMC_62 TSMC_110 TSMC_111 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW2 TSMC_91 TSMC_92 TSMC_112 TSMC_113 TSMC_101 VDDM VDDAI VSS TSMC_27 
+ TSMC_28 TSMC_59 TSMC_60 TSMC_114 TSMC_115 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW3 TSMC_89 TSMC_90 TSMC_116 TSMC_117 TSMC_101 VDDM VDDAI VSS TSMC_25 
+ TSMC_26 TSMC_57 TSMC_58 TSMC_118 TSMC_119 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW4 TSMC_87 TSMC_88 TSMC_120 TSMC_121 TSMC_101 VDDM VDDAI VSS TSMC_23 
+ TSMC_24 TSMC_55 TSMC_56 TSMC_122 TSMC_123 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW5 TSMC_85 TSMC_86 TSMC_124 TSMC_125 TSMC_101 VDDM VDDAI VSS TSMC_21 
+ TSMC_22 TSMC_53 TSMC_54 TSMC_126 TSMC_127 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW6 TSMC_83 TSMC_84 TSMC_128 TSMC_129 TSMC_101 VDDM VDDAI VSS TSMC_19 
+ TSMC_20 TSMC_51 TSMC_52 TSMC_130 TSMC_131 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW7 TSMC_81 TSMC_82 TSMC_132 TSMC_133 TSMC_101 VDDM VDDAI VSS TSMC_17 
+ TSMC_18 TSMC_49 TSMC_50 TSMC_134 TSMC_135 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW8 TSMC_79 TSMC_80 TSMC_136 TSMC_137 TSMC_101 VDDM VDDAI VSS TSMC_15 
+ TSMC_16 TSMC_47 TSMC_48 TSMC_138 TSMC_139 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW9 TSMC_77 TSMC_78 TSMC_140 TSMC_141 TSMC_101 VDDM VDDAI VSS TSMC_13 
+ TSMC_14 TSMC_45 TSMC_46 TSMC_142 TSMC_143 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW10 TSMC_75 TSMC_76 TSMC_144 TSMC_145 TSMC_101 VDDM VDDAI VSS TSMC_11 
+ TSMC_12 TSMC_43 TSMC_44 TSMC_146 TSMC_147 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW11 TSMC_73 TSMC_74 TSMC_148 TSMC_149 TSMC_101 VDDM VDDAI VSS TSMC_9 
+ TSMC_10 TSMC_41 TSMC_42 TSMC_150 TSMC_151 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW12 TSMC_71 TSMC_72 TSMC_152 TSMC_153 TSMC_101 VDDM VDDAI VSS TSMC_7 
+ TSMC_8 TSMC_39 TSMC_40 TSMC_154 TSMC_155 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW13 TSMC_69 TSMC_70 TSMC_156 TSMC_157 TSMC_101 VDDM VDDAI VSS TSMC_5 
+ TSMC_6 TSMC_37 TSMC_38 TSMC_158 TSMC_159 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW14 TSMC_67 TSMC_68 TSMC_160 TSMC_161 TSMC_101 VDDM VDDAI VSS TSMC_3 
+ TSMC_4 TSMC_35 TSMC_36 TSMC_162 TSMC_163 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROW15 TSMC_65 TSMC_66 TSMC_164 TSMC_165 TSMC_101 VDDM VDDAI VSS TSMC_1 
+ TSMC_2 TSMC_33 TSMC_34 TSMC_166 TSMC_167 VSS 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XTRKROWL TSMC_168 TSMC_169 TSMC_101 VDDM VDDAI VSS TSMC_102 TSMC_170 
+ TSMC_171 VSS S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X1 
XTRKROWR TSMC_97 TSMC_172 TSMC_101 VDDM VDDAI VSS TSMC_103 TSMC_173 
+ TSMC_174 VSS S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X1 
XTRKCTRL TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 
+ TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_100 TSMC_98 TSMC_99 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 
+ TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_101 VDDM VDDI VSS TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ S6ALLSVTFW8U20_RF_TRKCTRL 
.ENDS

.SUBCKT S6ALLSVTFW8U20_ARY4ROW TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 
+ TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 
+ TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 
+ TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 
+ TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 
+ TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 VDDM VDDAI VDDI VSS 
+ TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
XCOL0 TSMC_31 TSMC_32 TSMC_63 TSMC_64 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_95 TSMC_96 TSMC_127 TSMC_128 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL1 TSMC_29 TSMC_30 TSMC_61 TSMC_62 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_93 TSMC_94 TSMC_125 TSMC_126 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL2 TSMC_27 TSMC_28 TSMC_59 TSMC_60 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_91 TSMC_92 TSMC_123 TSMC_124 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL3 TSMC_25 TSMC_26 TSMC_57 TSMC_58 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_89 TSMC_90 TSMC_121 TSMC_122 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL4 TSMC_23 TSMC_24 TSMC_55 TSMC_56 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_87 TSMC_88 TSMC_119 TSMC_120 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL5 TSMC_21 TSMC_22 TSMC_53 TSMC_54 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_85 TSMC_86 TSMC_117 TSMC_118 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL6 TSMC_19 TSMC_20 TSMC_51 TSMC_52 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_83 TSMC_84 TSMC_115 TSMC_116 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL7 TSMC_17 TSMC_18 TSMC_49 TSMC_50 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_81 TSMC_82 TSMC_113 TSMC_114 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL8 TSMC_15 TSMC_16 TSMC_47 TSMC_48 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_79 TSMC_80 TSMC_111 TSMC_112 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL9 TSMC_13 TSMC_14 TSMC_45 TSMC_46 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_77 TSMC_78 TSMC_109 TSMC_110 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL10 TSMC_11 TSMC_12 TSMC_43 TSMC_44 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_75 TSMC_76 TSMC_107 TSMC_108 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL11 TSMC_9 TSMC_10 TSMC_41 TSMC_42 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_73 TSMC_74 TSMC_105 TSMC_106 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL12 TSMC_7 TSMC_8 TSMC_39 TSMC_40 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_71 TSMC_72 TSMC_103 TSMC_104 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL13 TSMC_5 TSMC_6 TSMC_37 TSMC_38 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_69 TSMC_70 TSMC_101 TSMC_102 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL14 TSMC_3 TSMC_4 TSMC_35 TSMC_36 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_67 TSMC_68 TSMC_99 TSMC_100 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL15 TSMC_1 TSMC_2 TSMC_33 TSMC_34 TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM 
+ VDDAI VSS TSMC_65 TSMC_66 TSMC_97 TSMC_98 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XTRKL TSMC_129 TSMC_192 TSMC_193 TSMC_180 TSMC_181 TSMC_130 TSMC_130 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM VDDAI VSS TSMC_176 TSMC_177 VSS 
+ TSMC_131 TSMC_188 TSMC_189 TSMC_190 TSMC_191 
+ S6ALLSVTFW8U20_D130_ARRAY_RBL_TRK_OFF_4X1 
XTRKR TSMC_132 TSMC_194 TSMC_195 TSMC_182 TSMC_183 TSMC_130 TSMC_130 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 VDDM VDDAI VSS TSMC_178 TSMC_179 VSS 
+ TSMC_133 TSMC_188 TSMC_189 TSMC_190 TSMC_191 
+ S6ALLSVTFW8U20_D130_ARRAY_RBL_TRK_OFF_4X1 
XDEC TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_134 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_187 TSMC_152 VDDM VDDI VDDI VSS TSMC_153 
+ TSMC_154 TSMC_155 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 
+ TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 TSMC_172 TSMC_173 TSMC_174 TSMC_175 
+ S6ALLSVTFW8U20_RF_XDEC4 
.ENDS

.SUBCKT S6ALLSVTFW8U20_ARY4ROW_TK TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 VDDM VDDAI 
+ VDDI VSS TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 
+ TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 
+ TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 
XCOL0 TSMC_31 TSMC_32 TSMC_63 TSMC_64 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_95 TSMC_96 TSMC_127 TSMC_128 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL1 TSMC_29 TSMC_30 TSMC_61 TSMC_62 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_93 TSMC_94 TSMC_125 TSMC_126 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL2 TSMC_27 TSMC_28 TSMC_59 TSMC_60 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_91 TSMC_92 TSMC_123 TSMC_124 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL3 TSMC_25 TSMC_26 TSMC_57 TSMC_58 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_89 TSMC_90 TSMC_121 TSMC_122 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL4 TSMC_23 TSMC_24 TSMC_55 TSMC_56 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_87 TSMC_88 TSMC_119 TSMC_120 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL5 TSMC_21 TSMC_22 TSMC_53 TSMC_54 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_85 TSMC_86 TSMC_117 TSMC_118 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL6 TSMC_19 TSMC_20 TSMC_51 TSMC_52 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_83 TSMC_84 TSMC_115 TSMC_116 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL7 TSMC_17 TSMC_18 TSMC_49 TSMC_50 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_81 TSMC_82 TSMC_113 TSMC_114 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL8 TSMC_15 TSMC_16 TSMC_47 TSMC_48 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_79 TSMC_80 TSMC_111 TSMC_112 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL9 TSMC_13 TSMC_14 TSMC_45 TSMC_46 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_77 TSMC_78 TSMC_109 TSMC_110 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL10 TSMC_11 TSMC_12 TSMC_43 TSMC_44 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_75 TSMC_76 TSMC_107 TSMC_108 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL11 TSMC_9 TSMC_10 TSMC_41 TSMC_42 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_73 TSMC_74 TSMC_105 TSMC_106 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL12 TSMC_7 TSMC_8 TSMC_39 TSMC_40 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_71 TSMC_72 TSMC_103 TSMC_104 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL13 TSMC_5 TSMC_6 TSMC_37 TSMC_38 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_69 TSMC_70 TSMC_101 TSMC_102 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL14 TSMC_3 TSMC_4 TSMC_35 TSMC_36 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_67 TSMC_68 TSMC_99 TSMC_100 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XCOL15 TSMC_1 TSMC_2 TSMC_33 TSMC_34 TSMC_186 TSMC_187 TSMC_188 TSMC_189 VDDM 
+ VDDAI VSS TSMC_65 TSMC_66 TSMC_97 TSMC_98 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_4X2 
XTRKL TSMC_129 TSMC_194 TSMC_195 TSMC_182 TSMC_183 TSMC_130 TSMC_130 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_180 TSMC_180 VDDM VDDAI VSS VSS 
+ TSMC_176 TSMC_177 TSMC_131 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_RBL_TRK_4X1 
XTRKR TSMC_196 TSMC_197 TSMC_198 TSMC_184 TSMC_185 TSMC_130 TSMC_130 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_181 TSMC_181 VDDM VDDAI VSS VSS 
+ TSMC_178 TSMC_179 TSMC_133 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 S6ALLSVTFW8U20_D130_ARRAY_RBL_TRK_4X1 
XDEC TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 
+ TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 
+ TSMC_214 TSMC_215 TSMC_134 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_152 VDDM VDDI VDDI VSS TSMC_153 
+ TSMC_154 TSMC_155 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 
+ TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_172 TSMC_173 TSMC_174 TSMC_175 
+ S6ALLSVTFW8U20_RF_XDEC4 
.ENDS

.SUBCKT S6ALLSVTFW8U20_LIO_LCTRL TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 
+ TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 
+ TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 
+ TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 VDDM VDDI VDDAI VSS 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 
+ TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 
+ TSMC_232 TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 
XLIO0 TSMC_31 TSMC_32 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_63 
+ TSMC_64 TSMC_95 TSMC_96 TSMC_213 VDDM VDDAI VDDI VSS TSMC_127 
+ TSMC_128 TSMC_159 TSMC_160 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO1 TSMC_29 TSMC_30 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_61 
+ TSMC_62 TSMC_93 TSMC_94 TSMC_213 VDDM VDDAI VDDI VSS TSMC_125 
+ TSMC_126 TSMC_157 TSMC_158 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO2 TSMC_27 TSMC_28 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_59 
+ TSMC_60 TSMC_91 TSMC_92 TSMC_213 VDDM VDDAI VDDI VSS TSMC_123 
+ TSMC_124 TSMC_155 TSMC_156 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO3 TSMC_25 TSMC_26 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_57 
+ TSMC_58 TSMC_89 TSMC_90 TSMC_213 VDDM VDDAI VDDI VSS TSMC_121 
+ TSMC_122 TSMC_153 TSMC_154 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO4 TSMC_23 TSMC_24 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_55 
+ TSMC_56 TSMC_87 TSMC_88 TSMC_213 VDDM VDDAI VDDI VSS TSMC_119 
+ TSMC_120 TSMC_151 TSMC_152 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO5 TSMC_21 TSMC_22 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_53 
+ TSMC_54 TSMC_85 TSMC_86 TSMC_213 VDDM VDDAI VDDI VSS TSMC_117 
+ TSMC_118 TSMC_149 TSMC_150 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO6 TSMC_19 TSMC_20 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_51 
+ TSMC_52 TSMC_83 TSMC_84 TSMC_213 VDDM VDDAI VDDI VSS TSMC_115 
+ TSMC_116 TSMC_147 TSMC_148 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO7 TSMC_17 TSMC_18 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_49 
+ TSMC_50 TSMC_81 TSMC_82 TSMC_213 VDDM VDDAI VDDI VSS TSMC_113 
+ TSMC_114 TSMC_145 TSMC_146 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO8 TSMC_15 TSMC_16 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_47 
+ TSMC_48 TSMC_79 TSMC_80 TSMC_213 VDDM VDDAI VDDI VSS TSMC_111 
+ TSMC_112 TSMC_143 TSMC_144 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO9 TSMC_13 TSMC_14 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_45 
+ TSMC_46 TSMC_77 TSMC_78 TSMC_213 VDDM VDDAI VDDI VSS TSMC_109 
+ TSMC_110 TSMC_141 TSMC_142 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO10 TSMC_11 TSMC_12 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_43 TSMC_44 TSMC_75 TSMC_76 TSMC_213 VDDM VDDAI VDDI VSS TSMC_107 
+ TSMC_108 TSMC_139 TSMC_140 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO11 TSMC_9 TSMC_10 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_41 TSMC_42 TSMC_73 TSMC_74 TSMC_213 VDDM VDDAI VDDI VSS TSMC_105 
+ TSMC_106 TSMC_137 TSMC_138 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO12 TSMC_7 TSMC_8 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_39 TSMC_40 TSMC_71 TSMC_72 TSMC_213 VDDM VDDAI VDDI VSS TSMC_103 
+ TSMC_104 TSMC_135 TSMC_136 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO13 TSMC_5 TSMC_6 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_37 TSMC_38 TSMC_69 TSMC_70 TSMC_213 VDDM VDDAI VDDI VSS TSMC_101 
+ TSMC_102 TSMC_133 TSMC_134 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO14 TSMC_3 TSMC_4 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_35 TSMC_36 TSMC_67 TSMC_68 TSMC_213 VDDM VDDAI VDDI VSS TSMC_99 
+ TSMC_100 TSMC_131 TSMC_132 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XLIO15 TSMC_1 TSMC_2 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_33 TSMC_34 TSMC_65 TSMC_66 TSMC_213 VDDM VDDAI VDDI VSS TSMC_97 
+ TSMC_98 TSMC_129 TSMC_130 S6ALLSVTFW8U20_RF_LIOX2_72_V1 
XTROLIOL TSMC_239 TSMC_161 TSMC_237 TSMC_162 TSMC_163 TSMC_242 TSMC_243 
+ TSMC_244 TSMC_247 TSMC_248 TSMC_249 TSMC_245 TSMC_246 TSMC_164 
+ TSMC_165 TSMC_241 TSMC_167 TSMC_213 VDDM VDDAI VDDI VSS TSMC_250 
+ TSMC_169 TSMC_251 TSMC_171 TSMC_172 TSMC_173 
+ S6ALLSVTFW8U20_RF_TRKLIOX2_72_V1 
XTROLIOR TSMC_239 TSMC_174 TSMC_252 TSMC_175 TSMC_176 TSMC_242 TSMC_243 
+ TSMC_244 TSMC_247 TSMC_248 TSMC_249 TSMC_245 TSMC_246 TSMC_164 
+ TSMC_165 TSMC_241 TSMC_177 TSMC_213 VDDM VDDAI VDDI VSS TSMC_178 
+ TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ S6ALLSVTFW8U20_RF_TRKLIOX2_72_V1 
XLCTRL TSMC_238 TSMC_184 TSMC_185 TSMC_239 TSMC_240 TSMC_253 TSMC_254 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_247 TSMC_248 TSMC_249 TSMC_186 TSMC_187 
+ TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_245 TSMC_246 TSMC_164 
+ TSMC_255 TSMC_192 TSMC_166 TSMC_193 TSMC_194 TSMC_195 TSMC_196 
+ TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 
+ TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_213 TSMC_165 TSMC_214 TSMC_215 VDDM VDDI VSS TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 
+ TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 
+ TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 TSMC_236 
+ S6ALLSVTFW8U20_RF_LCTRL 
.ENDS

.SUBCKT S6ALLSVTFW8U20_WRITE_TRAKING TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 VDDM VDDI VDDAI VSS TSMC_140 TSMC_141 TSMC_142 TSMC_143 
+ TSMC_144 
XRWLLD0 TSMC_31 TSMC_32 TSMC_63 TSMC_64 VSS VDDM VDDAI VSS TSMC_127 TSMC_128 
+ TSMC_95 TSMC_96 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD1 TSMC_29 TSMC_30 TSMC_61 TSMC_62 VSS VDDM VDDAI VSS TSMC_125 TSMC_126 
+ TSMC_93 TSMC_94 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD2 TSMC_27 TSMC_28 TSMC_59 TSMC_60 VSS VDDM VDDAI VSS TSMC_123 TSMC_124 
+ TSMC_91 TSMC_92 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD3 TSMC_25 TSMC_26 TSMC_57 TSMC_58 VSS VDDM VDDAI VSS TSMC_121 TSMC_122 
+ TSMC_89 TSMC_90 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD4 TSMC_23 TSMC_24 TSMC_55 TSMC_56 VSS VDDM VDDAI VSS TSMC_119 TSMC_120 
+ TSMC_87 TSMC_88 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD5 TSMC_21 TSMC_22 TSMC_53 TSMC_54 VSS VDDM VDDAI VSS TSMC_117 
+ TSMC_118 TSMC_85 TSMC_86 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD6 TSMC_19 TSMC_20 TSMC_51 TSMC_52 VSS VDDM VDDAI VSS TSMC_115 
+ TSMC_116 TSMC_83 TSMC_84 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD7 TSMC_17 TSMC_18 TSMC_49 TSMC_50 VSS VDDM VDDAI VSS TSMC_113 
+ TSMC_114 TSMC_81 TSMC_82 TSMC_145 TSMC_146 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD8 TSMC_15 TSMC_16 TSMC_47 TSMC_48 VSS VDDM VDDAI VSS TSMC_111 
+ TSMC_112 TSMC_79 TSMC_80 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD9 TSMC_13 TSMC_14 TSMC_45 TSMC_46 VSS VDDM VDDAI VSS TSMC_109 
+ TSMC_110 TSMC_77 TSMC_78 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD10 TSMC_11 TSMC_12 TSMC_43 TSMC_44 VSS VDDM VDDAI VSS TSMC_107 
+ TSMC_108 TSMC_75 TSMC_76 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD11 TSMC_9 TSMC_10 TSMC_41 TSMC_42 VSS VDDM VDDAI VSS TSMC_105 
+ TSMC_106 TSMC_73 TSMC_74 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD12 TSMC_7 TSMC_8 TSMC_39 TSMC_40 VSS VDDM VDDAI VSS TSMC_103 
+ TSMC_104 TSMC_71 TSMC_72 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD13 TSMC_5 TSMC_6 TSMC_37 TSMC_38 VSS VDDM VDDAI VSS TSMC_101 
+ TSMC_102 TSMC_69 TSMC_70 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD14 TSMC_3 TSMC_4 TSMC_35 TSMC_36 VSS VDDM VDDAI VSS TSMC_99 
+ TSMC_100 TSMC_67 TSMC_68 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLD15 TSMC_1 TSMC_2 TSMC_33 TSMC_34 VSS VDDM VDDAI VSS TSMC_97 
+ TSMC_98 TSMC_65 TSMC_66 TSMC_148 TSMC_149 TSMC_147 
+ S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X2 
XRWLLDL TSMC_129 TSMC_130 VSS VDDM VDDAI VSS TSMC_150 TSMC_131 TSMC_151 
+ TSMC_147 S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X1 
XRWLLDR TSMC_133 TSMC_130 VSS VDDM VDDAI VSS TSMC_152 TSMC_134 TSMC_151 
+ TSMC_147 S6ALLSVTFW8U20_D130_ARRAY_RWL_TRK_X1 
XDECCAP TSMC_153 TSMC_139 TSMC_136 TSMC_137 TSMC_138 VDDM VDDI VSS TSMC_131 
+ TSMC_135 TSMC_132 TSMC_140 TSMC_147 TSMC_147 
+ S6ALLSVTFW8U20_RF_XDECCAP 
.ENDS

.SUBCKT TS6N16FFCLLSVTA8X32M1FW D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] 
+ D[23] D[22] D[21] D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] 
+ D[10] D[9] D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] Q[31] Q[30] Q[29] 
+ Q[28] Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] Q[16] 
+ Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] 
+ Q[1] Q[0] BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] BWEB[25] 
+ BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] BWEB[18] BWEB[17] 
+ BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] BWEB[11] BWEB[10] BWEB[9] 
+ BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] BWEB[3] BWEB[2] BWEB[1] BWEB[0] AB[2] 
+ AB[1] AB[0] CLKR REB AA[2] AA[1] AA[0] CLKW WEB KP[2] KP[1] KP[0] WCT[1] 
+ WCT[0] RCT[1] RCT[0] VDD VSS 
XPIN_ROW D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] D[22] D[21] 
+ D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] D[10] D[9] 
+ D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] Q[31] Q[30] Q[29] Q[28] 
+ Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] Q[16] 
+ Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] 
+ Q[2] Q[1] Q[0] BWEB[31] BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] 
+ BWEB[25] BWEB[24] BWEB[23] BWEB[22] BWEB[21] BWEB[20] BWEB[19] 
+ BWEB[18] BWEB[17] BWEB[16] BWEB[15] BWEB[14] BWEB[13] BWEB[12] 
+ BWEB[11] BWEB[10] BWEB[9] BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] 
+ BWEB[3] BWEB[2] BWEB[1] BWEB[0] TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 AB[2] AB[1] AB[0] CLKR REB TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 AA[2] AA[1] AA[0] CLKW WEB KP[2] KP[1] 
+ KP[0] TSMC_1 TSMC_2 TSMC_1 RCT[1] RCT[0] WCT[1] WCT[0] TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 VSS TSMC_3 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_2 TSMC_2 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_4 
+ TSMC_5 TSMC_6 S6ALLSVTFW8U20_PIN_ROW 
XGCTRL_GIO CLKR CLKW D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] 
+ D[22] D[21] D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] 
+ D[10] D[9] D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 KP[2] KP[1] KP[0] 
+ TSMC_72 TSMC_73 TSMC_74 TSMC_1 TSMC_2 TSMC_1 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_1 Q[31] Q[30] Q[29] Q[28] Q[27] Q[26] Q[25] Q[24] 
+ Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17] Q[16] Q[15] Q[14] Q[13] Q[12] 
+ Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] RCT[1] 
+ RCT[0] REB TSMC_80 TSMC_1 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
+ TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 AB[2] AB[1] AB[0] TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_2 TSMC_1 TSMC_100 VDD VDD VSS TSMC_101 TSMC_102 TSMC_103 
+ TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 
+ TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 
+ TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 WCT[1] WCT[0] WEB BWEB[31] BWEB[30] 
+ BWEB[29] BWEB[28] BWEB[27] BWEB[26] BWEB[25] BWEB[24] BWEB[23] 
+ BWEB[22] BWEB[21] BWEB[20] BWEB[19] BWEB[18] BWEB[17] BWEB[16] 
+ BWEB[15] BWEB[14] BWEB[13] BWEB[12] BWEB[11] BWEB[10] BWEB[9] 
+ BWEB[8] BWEB[7] BWEB[6] BWEB[5] BWEB[4] BWEB[3] BWEB[2] BWEB[1] 
+ BWEB[0] TSMC_165 TSMC_1 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_171 
+ TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 
+ TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 AA[2] AA[1] AA[0] TSMC_1 TSMC_1 TSMC_1 TSMC_185 
+ TSMC_1 TSMC_3 TSMC_186 TSMC_2 TSMC_187 TSMC_2 TSMC_2 VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_1 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 
+ TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_2 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 
+ TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 
+ TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_1 S6ALLSVTFW8U20_GCTRL_GIO 
XROW_TRACKING TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_101 TSMC_102 TSMC_103 
+ TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 VDD 
+ VDD VDD VSS TSMC_80 TSMC_80 TSMC_1 TSMC_100 TSMC_252 TSMC_253 
+ S6ALLSVTFW8U20_ROW_TRACKING 
XARY4ROW_SEG0_ARY0 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 
+ TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 
+ TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_286 
+ TSMC_287 TSMC_78 TSMC_71 TSMC_288 TSMC_289 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_1 TSMC_1 VDD VDD VDD VSS 
+ TSMC_165 TSMC_166 TSMC_290 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_91 TSMC_95 TSMC_176 
+ TSMC_180 TSMC_252 TSMC_291 TSMC_253 TSMC_292 TSMC_293 
+ TSMC_294 TSMC_295 TSMC_296 S6ALLSVTFW8U20_ARY4ROW 
XARY4ROW_TK_SEG0_ARY1 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 
+ TSMC_70 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 
+ TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 
+ TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 
+ TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 
+ TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 
+ TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_286 
+ TSMC_287 TSMC_78 TSMC_71 TSMC_288 TSMC_289 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_1 TSMC_1 VDD VDD VDD VSS 
+ TSMC_165 TSMC_166 TSMC_290 TSMC_169 TSMC_170 TSMC_171 TSMC_172 
+ TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 
+ TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_90 TSMC_95 TSMC_175 
+ TSMC_180 TSMC_291 TSMC_297 TSMC_292 TSMC_298 TSMC_100 
+ TSMC_100 TSMC_294 TSMC_299 TSMC_296 TSMC_300 
+ S6ALLSVTFW8U20_ARY4ROW_TK 
XLIO_LCTRL_SEG0 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 
+ TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 
+ TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 
+ TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 
+ TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 TSMC_306 TSMC_307 
+ TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 TSMC_313 
+ TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 
+ TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_133 
+ TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 
+ TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 
+ TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 TSMC_155 
+ TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 
+ TSMC_163 TSMC_164 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 
+ TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 
+ TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_333 TSMC_286 
+ TSMC_333 TSMC_1 TSMC_287 TSMC_80 TSMC_100 TSMC_1 TSMC_1 TSMC_1 
+ TSMC_78 TSMC_79 TSMC_100 TSMC_334 TSMC_71 TSMC_334 TSMC_100 TSMC_1 
+ TSMC_1 TSMC_1 VDD TSMC_185 TSMC_100 TSMC_95 TSMC_95 TSMC_72 TSMC_73 TSMC_74 
+ TSMC_75 TSMC_76 TSMC_77 TSMC_1 TSMC_335 TSMC_81 TSMC_289 TSMC_84 
+ TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 
+ TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_1 TSMC_1 
+ TSMC_94 TSMC_94 VDD VDD VDD VSS TSMC_165 TSMC_166 TSMC_290 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_80 TSMC_165 TSMC_336 TSMC_187 TSMC_1 TSMC_337 TSMC_80 
+ S6ALLSVTFW8U20_LIO_LCTRL 
XWRITE_TRAKING TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 
+ TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 
+ TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 
+ TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 
+ TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_101 
+ TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 
+ TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 TSMC_115 
+ TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 
+ TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_286 
+ TSMC_287 TSMC_78 TSMC_79 TSMC_71 TSMC_288 TSMC_185 TSMC_80 TSMC_335 TSMC_1 
+ TSMC_1 VDD VDD VDD VSS TSMC_165 TSMC_297 TSMC_298 TSMC_299 
+ TSMC_300 S6ALLSVTFW8U20_WRITE_TRAKING 
.ENDS


