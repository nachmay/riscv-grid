# Created by MC2 : Version 2013.12.00.f on 2025/06/22, 17:57:14

#*********************************************************************************************************************/
# Technology     : TSMC 16nm CMOS Logic FinFet Compact (FFC) Low Leakage HKMG                          */
# Memory Type    : TSMC 16nm FFC Single Port SRAM with d0907 bit cell                     */
# Library Name   : ts1n16ffcllsvta1024x32m4sw (user specify : ts1n16ffcllsvta1024x32m4sw)            */
# Library Version: 120a                                                */
# Generated Time : 2025/06/22, 17:57:08                                        */
#*********************************************************************************************************************/
#                                                            */
# STATEMENT OF USE                                                    */
#                                                            */
# This information contains confidential and proprietary information of TSMC.                    */
# No part of this information may be reproduced, transmitted, transcribed,                        */
# stored in a retrieval system, or translated into any human or computer                        */
# language, in any form or by any means, electronic, mechanical, magnetic,                        */
# optical, chemical, manual, or otherwise, without the prior written permission                    */
# of TSMC. This information was prepared for informational purpose and is for                    */
# use by TSMC's customers only. TSMC reserves the right to make changes in the                    */
# information at any time and without notice.                                    */
#                                                            */
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N16FFCLLSVTA1024X32M4SW
	CLASS BLOCK ;
	FOREIGN TS1N16FFCLLSVTA1024X32M4SW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 60.575 BY 79.344 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 34.952 60.575 35.032 ;
			LAYER M2 ;
			RECT 60.327 34.952 60.575 35.032 ;
			LAYER M3 ;
			RECT 60.327 34.952 60.575 35.032 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 33.608 60.575 33.688 ;
			LAYER M2 ;
			RECT 60.327 33.608 60.575 33.688 ;
			LAYER M3 ;
			RECT 60.327 33.608 60.575 33.688 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 43.976 60.575 44.056 ;
			LAYER M2 ;
			RECT 60.327 43.976 60.575 44.056 ;
			LAYER M3 ;
			RECT 60.327 43.976 60.575 44.056 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 43.208 60.575 43.288 ;
			LAYER M2 ;
			RECT 60.327 43.208 60.575 43.288 ;
			LAYER M3 ;
			RECT 60.327 43.208 60.575 43.288 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 42.632 60.575 42.712 ;
			LAYER M2 ;
			RECT 60.327 42.632 60.575 42.712 ;
			LAYER M3 ;
			RECT 60.327 42.632 60.575 42.712 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 39.944 60.575 40.024 ;
			LAYER M2 ;
			RECT 60.327 39.944 60.575 40.024 ;
			LAYER M3 ;
			RECT 60.327 39.944 60.575 40.024 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 40.712 60.575 40.792 ;
			LAYER M2 ;
			RECT 60.327 40.712 60.575 40.792 ;
			LAYER M3 ;
			RECT 60.327 40.712 60.575 40.792 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 41.864 60.575 41.944 ;
			LAYER M2 ;
			RECT 60.327 41.864 60.575 41.944 ;
			LAYER M3 ;
			RECT 60.327 41.864 60.575 41.944 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 36.488 60.575 36.568 ;
			LAYER M2 ;
			RECT 60.327 36.488 60.575 36.568 ;
			LAYER M3 ;
			RECT 60.327 36.488 60.575 36.568 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 35.144 60.575 35.224 ;
			LAYER M2 ;
			RECT 60.327 35.144 60.575 35.224 ;
			LAYER M3 ;
			RECT 60.327 35.144 60.575 35.224 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.834200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.362400 LAYER M2 ;
		ANTENNAMAXAREACAR 11.423200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.199400 LAYER M3 ;
		ANTENNAMAXAREACAR 33.069400 LAYER M3 ;
	END A[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 1.976 60.575 2.056 ;
			LAYER M2 ;
			RECT 60.327 1.976 60.575 2.056 ;
			LAYER M3 ;
			RECT 60.327 1.976 60.575 2.056 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 3.992 60.575 4.072 ;
			LAYER M2 ;
			RECT 60.327 3.992 60.575 4.072 ;
			LAYER M3 ;
			RECT 60.327 3.992 60.575 4.072 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 6.008 60.575 6.088 ;
			LAYER M2 ;
			RECT 60.327 6.008 60.575 6.088 ;
			LAYER M3 ;
			RECT 60.327 6.008 60.575 6.088 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 8.024 60.575 8.104 ;
			LAYER M2 ;
			RECT 60.327 8.024 60.575 8.104 ;
			LAYER M3 ;
			RECT 60.327 8.024 60.575 8.104 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 10.040 60.575 10.120 ;
			LAYER M2 ;
			RECT 60.327 10.040 60.575 10.120 ;
			LAYER M3 ;
			RECT 60.327 10.040 60.575 10.120 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 12.056 60.575 12.136 ;
			LAYER M2 ;
			RECT 60.327 12.056 60.575 12.136 ;
			LAYER M3 ;
			RECT 60.327 12.056 60.575 12.136 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 14.072 60.575 14.152 ;
			LAYER M2 ;
			RECT 60.327 14.072 60.575 14.152 ;
			LAYER M3 ;
			RECT 60.327 14.072 60.575 14.152 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 16.088 60.575 16.168 ;
			LAYER M2 ;
			RECT 60.327 16.088 60.575 16.168 ;
			LAYER M3 ;
			RECT 60.327 16.088 60.575 16.168 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 18.104 60.575 18.184 ;
			LAYER M2 ;
			RECT 60.327 18.104 60.575 18.184 ;
			LAYER M3 ;
			RECT 60.327 18.104 60.575 18.184 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 20.120 60.575 20.200 ;
			LAYER M2 ;
			RECT 60.327 20.120 60.575 20.200 ;
			LAYER M3 ;
			RECT 60.327 20.120 60.575 20.200 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 22.136 60.575 22.216 ;
			LAYER M2 ;
			RECT 60.327 22.136 60.575 22.216 ;
			LAYER M3 ;
			RECT 60.327 22.136 60.575 22.216 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 24.152 60.575 24.232 ;
			LAYER M2 ;
			RECT 60.327 24.152 60.575 24.232 ;
			LAYER M3 ;
			RECT 60.327 24.152 60.575 24.232 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 26.168 60.575 26.248 ;
			LAYER M2 ;
			RECT 60.327 26.168 60.575 26.248 ;
			LAYER M3 ;
			RECT 60.327 26.168 60.575 26.248 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 28.184 60.575 28.264 ;
			LAYER M2 ;
			RECT 60.327 28.184 60.575 28.264 ;
			LAYER M3 ;
			RECT 60.327 28.184 60.575 28.264 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 30.200 60.575 30.280 ;
			LAYER M2 ;
			RECT 60.327 30.200 60.575 30.280 ;
			LAYER M3 ;
			RECT 60.327 30.200 60.575 30.280 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 32.216 60.575 32.296 ;
			LAYER M2 ;
			RECT 60.327 32.216 60.575 32.296 ;
			LAYER M3 ;
			RECT 60.327 32.216 60.575 32.296 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 47.096 60.575 47.176 ;
			LAYER M2 ;
			RECT 60.327 47.096 60.575 47.176 ;
			LAYER M3 ;
			RECT 60.327 47.096 60.575 47.176 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 49.112 60.575 49.192 ;
			LAYER M2 ;
			RECT 60.327 49.112 60.575 49.192 ;
			LAYER M3 ;
			RECT 60.327 49.112 60.575 49.192 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 51.128 60.575 51.208 ;
			LAYER M2 ;
			RECT 60.327 51.128 60.575 51.208 ;
			LAYER M3 ;
			RECT 60.327 51.128 60.575 51.208 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 53.144 60.575 53.224 ;
			LAYER M2 ;
			RECT 60.327 53.144 60.575 53.224 ;
			LAYER M3 ;
			RECT 60.327 53.144 60.575 53.224 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 55.160 60.575 55.240 ;
			LAYER M2 ;
			RECT 60.327 55.160 60.575 55.240 ;
			LAYER M3 ;
			RECT 60.327 55.160 60.575 55.240 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 57.176 60.575 57.256 ;
			LAYER M2 ;
			RECT 60.327 57.176 60.575 57.256 ;
			LAYER M3 ;
			RECT 60.327 57.176 60.575 57.256 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 59.192 60.575 59.272 ;
			LAYER M2 ;
			RECT 60.327 59.192 60.575 59.272 ;
			LAYER M3 ;
			RECT 60.327 59.192 60.575 59.272 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 61.208 60.575 61.288 ;
			LAYER M2 ;
			RECT 60.327 61.208 60.575 61.288 ;
			LAYER M3 ;
			RECT 60.327 61.208 60.575 61.288 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 63.224 60.575 63.304 ;
			LAYER M2 ;
			RECT 60.327 63.224 60.575 63.304 ;
			LAYER M3 ;
			RECT 60.327 63.224 60.575 63.304 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 65.240 60.575 65.320 ;
			LAYER M2 ;
			RECT 60.327 65.240 60.575 65.320 ;
			LAYER M3 ;
			RECT 60.327 65.240 60.575 65.320 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 67.256 60.575 67.336 ;
			LAYER M2 ;
			RECT 60.327 67.256 60.575 67.336 ;
			LAYER M3 ;
			RECT 60.327 67.256 60.575 67.336 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 69.272 60.575 69.352 ;
			LAYER M2 ;
			RECT 60.327 69.272 60.575 69.352 ;
			LAYER M3 ;
			RECT 60.327 69.272 60.575 69.352 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 71.288 60.575 71.368 ;
			LAYER M2 ;
			RECT 60.327 71.288 60.575 71.368 ;
			LAYER M3 ;
			RECT 60.327 71.288 60.575 71.368 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 73.304 60.575 73.384 ;
			LAYER M2 ;
			RECT 60.327 73.304 60.575 73.384 ;
			LAYER M3 ;
			RECT 60.327 73.304 60.575 73.384 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 75.320 60.575 75.400 ;
			LAYER M2 ;
			RECT 60.327 75.320 60.575 75.400 ;
			LAYER M3 ;
			RECT 60.327 75.320 60.575 75.400 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 77.336 60.575 77.416 ;
			LAYER M2 ;
			RECT 60.327 77.336 60.575 77.416 ;
			LAYER M3 ;
			RECT 60.327 77.336 60.575 77.416 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.093800 LAYER M1 ;
		ANTENNAMAXAREACAR 9.051800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.215000 LAYER M3 ;
		ANTENNAMAXAREACAR 128.793000 LAYER M3 ;
	END BWEB[31]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 36.680 60.575 36.760 ;
			LAYER M2 ;
			RECT 60.327 36.680 60.575 36.760 ;
			LAYER M3 ;
			RECT 60.327 36.680 60.575 36.760 ;
		END
		ANTENNAGATEAREA 0.010000 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081400 LAYER M1 ;
		ANTENNAMAXAREACAR 2.270000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.204800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010000 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127600 LAYER M2 ;
		ANTENNAMAXAREACAR 9.590000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.409600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010000 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.158200 LAYER M3 ;
		ANTENNAMAXAREACAR 25.420000 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 38.984 60.575 39.064 ;
			LAYER M2 ;
			RECT 60.327 38.984 60.575 39.064 ;
			LAYER M3 ;
			RECT 60.327 38.984 60.575 39.064 ;
		END
		ANTENNAGATEAREA 0.284200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 2.071400 LAYER M1 ;
		ANTENNAMAXAREACAR 12.657200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.061400 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.284200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 3.218800 LAYER M2 ;
		ANTENNAMAXAREACAR 73.469000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.031800 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.789800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.284200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.817000 LAYER M3 ;
		ANTENNAMAXAREACAR 83.379800 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 2.360 60.575 2.440 ;
			LAYER M2 ;
			RECT 60.327 2.360 60.575 2.440 ;
			LAYER M3 ;
			RECT 60.327 2.360 60.575 2.440 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 4.376 60.575 4.456 ;
			LAYER M2 ;
			RECT 60.327 4.376 60.575 4.456 ;
			LAYER M3 ;
			RECT 60.327 4.376 60.575 4.456 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 6.392 60.575 6.472 ;
			LAYER M2 ;
			RECT 60.327 6.392 60.575 6.472 ;
			LAYER M3 ;
			RECT 60.327 6.392 60.575 6.472 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 8.408 60.575 8.488 ;
			LAYER M2 ;
			RECT 60.327 8.408 60.575 8.488 ;
			LAYER M3 ;
			RECT 60.327 8.408 60.575 8.488 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 10.424 60.575 10.504 ;
			LAYER M2 ;
			RECT 60.327 10.424 60.575 10.504 ;
			LAYER M3 ;
			RECT 60.327 10.424 60.575 10.504 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 12.440 60.575 12.520 ;
			LAYER M2 ;
			RECT 60.327 12.440 60.575 12.520 ;
			LAYER M3 ;
			RECT 60.327 12.440 60.575 12.520 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 14.456 60.575 14.536 ;
			LAYER M2 ;
			RECT 60.327 14.456 60.575 14.536 ;
			LAYER M3 ;
			RECT 60.327 14.456 60.575 14.536 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 16.472 60.575 16.552 ;
			LAYER M2 ;
			RECT 60.327 16.472 60.575 16.552 ;
			LAYER M3 ;
			RECT 60.327 16.472 60.575 16.552 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 18.488 60.575 18.568 ;
			LAYER M2 ;
			RECT 60.327 18.488 60.575 18.568 ;
			LAYER M3 ;
			RECT 60.327 18.488 60.575 18.568 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 20.504 60.575 20.584 ;
			LAYER M2 ;
			RECT 60.327 20.504 60.575 20.584 ;
			LAYER M3 ;
			RECT 60.327 20.504 60.575 20.584 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 22.520 60.575 22.600 ;
			LAYER M2 ;
			RECT 60.327 22.520 60.575 22.600 ;
			LAYER M3 ;
			RECT 60.327 22.520 60.575 22.600 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 24.536 60.575 24.616 ;
			LAYER M2 ;
			RECT 60.327 24.536 60.575 24.616 ;
			LAYER M3 ;
			RECT 60.327 24.536 60.575 24.616 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 26.552 60.575 26.632 ;
			LAYER M2 ;
			RECT 60.327 26.552 60.575 26.632 ;
			LAYER M3 ;
			RECT 60.327 26.552 60.575 26.632 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 28.568 60.575 28.648 ;
			LAYER M2 ;
			RECT 60.327 28.568 60.575 28.648 ;
			LAYER M3 ;
			RECT 60.327 28.568 60.575 28.648 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 30.584 60.575 30.664 ;
			LAYER M2 ;
			RECT 60.327 30.584 60.575 30.664 ;
			LAYER M3 ;
			RECT 60.327 30.584 60.575 30.664 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 32.600 60.575 32.680 ;
			LAYER M2 ;
			RECT 60.327 32.600 60.575 32.680 ;
			LAYER M3 ;
			RECT 60.327 32.600 60.575 32.680 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 47.480 60.575 47.560 ;
			LAYER M2 ;
			RECT 60.327 47.480 60.575 47.560 ;
			LAYER M3 ;
			RECT 60.327 47.480 60.575 47.560 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 49.496 60.575 49.576 ;
			LAYER M2 ;
			RECT 60.327 49.496 60.575 49.576 ;
			LAYER M3 ;
			RECT 60.327 49.496 60.575 49.576 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 51.512 60.575 51.592 ;
			LAYER M2 ;
			RECT 60.327 51.512 60.575 51.592 ;
			LAYER M3 ;
			RECT 60.327 51.512 60.575 51.592 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 53.528 60.575 53.608 ;
			LAYER M2 ;
			RECT 60.327 53.528 60.575 53.608 ;
			LAYER M3 ;
			RECT 60.327 53.528 60.575 53.608 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 55.544 60.575 55.624 ;
			LAYER M2 ;
			RECT 60.327 55.544 60.575 55.624 ;
			LAYER M3 ;
			RECT 60.327 55.544 60.575 55.624 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 57.560 60.575 57.640 ;
			LAYER M2 ;
			RECT 60.327 57.560 60.575 57.640 ;
			LAYER M3 ;
			RECT 60.327 57.560 60.575 57.640 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 59.576 60.575 59.656 ;
			LAYER M2 ;
			RECT 60.327 59.576 60.575 59.656 ;
			LAYER M3 ;
			RECT 60.327 59.576 60.575 59.656 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 61.592 60.575 61.672 ;
			LAYER M2 ;
			RECT 60.327 61.592 60.575 61.672 ;
			LAYER M3 ;
			RECT 60.327 61.592 60.575 61.672 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 63.608 60.575 63.688 ;
			LAYER M2 ;
			RECT 60.327 63.608 60.575 63.688 ;
			LAYER M3 ;
			RECT 60.327 63.608 60.575 63.688 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 65.624 60.575 65.704 ;
			LAYER M2 ;
			RECT 60.327 65.624 60.575 65.704 ;
			LAYER M3 ;
			RECT 60.327 65.624 60.575 65.704 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 67.640 60.575 67.720 ;
			LAYER M2 ;
			RECT 60.327 67.640 60.575 67.720 ;
			LAYER M3 ;
			RECT 60.327 67.640 60.575 67.720 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 69.656 60.575 69.736 ;
			LAYER M2 ;
			RECT 60.327 69.656 60.575 69.736 ;
			LAYER M3 ;
			RECT 60.327 69.656 60.575 69.736 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 71.672 60.575 71.752 ;
			LAYER M2 ;
			RECT 60.327 71.672 60.575 71.752 ;
			LAYER M3 ;
			RECT 60.327 71.672 60.575 71.752 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 73.688 60.575 73.768 ;
			LAYER M2 ;
			RECT 60.327 73.688 60.575 73.768 ;
			LAYER M3 ;
			RECT 60.327 73.688 60.575 73.768 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 75.704 60.575 75.784 ;
			LAYER M2 ;
			RECT 60.327 75.704 60.575 75.784 ;
			LAYER M3 ;
			RECT 60.327 75.704 60.575 75.784 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 77.720 60.575 77.800 ;
			LAYER M2 ;
			RECT 60.327 77.720 60.575 77.800 ;
			LAYER M3 ;
			RECT 60.327 77.720 60.575 77.800 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.111400 LAYER M1 ;
		ANTENNAMAXAREACAR 16.638000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.882800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.127400 LAYER M2 ;
		ANTENNAMAXAREACAR 40.517200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.765600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.232000 LAYER M3 ;
		ANTENNAMAXAREACAR 126.955000 LAYER M3 ;
	END D[31]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 1.208 60.575 1.288 ;
			LAYER M2 ;
			RECT 60.327 1.208 60.575 1.288 ;
			LAYER M3 ;
			RECT 60.327 1.208 60.575 1.288 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 3.224 60.575 3.304 ;
			LAYER M2 ;
			RECT 60.327 3.224 60.575 3.304 ;
			LAYER M3 ;
			RECT 60.327 3.224 60.575 3.304 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 5.240 60.575 5.320 ;
			LAYER M2 ;
			RECT 60.327 5.240 60.575 5.320 ;
			LAYER M3 ;
			RECT 60.327 5.240 60.575 5.320 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 7.256 60.575 7.336 ;
			LAYER M2 ;
			RECT 60.327 7.256 60.575 7.336 ;
			LAYER M3 ;
			RECT 60.327 7.256 60.575 7.336 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 9.272 60.575 9.352 ;
			LAYER M2 ;
			RECT 60.327 9.272 60.575 9.352 ;
			LAYER M3 ;
			RECT 60.327 9.272 60.575 9.352 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 11.288 60.575 11.368 ;
			LAYER M2 ;
			RECT 60.327 11.288 60.575 11.368 ;
			LAYER M3 ;
			RECT 60.327 11.288 60.575 11.368 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 13.304 60.575 13.384 ;
			LAYER M2 ;
			RECT 60.327 13.304 60.575 13.384 ;
			LAYER M3 ;
			RECT 60.327 13.304 60.575 13.384 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 15.320 60.575 15.400 ;
			LAYER M2 ;
			RECT 60.327 15.320 60.575 15.400 ;
			LAYER M3 ;
			RECT 60.327 15.320 60.575 15.400 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 17.336 60.575 17.416 ;
			LAYER M2 ;
			RECT 60.327 17.336 60.575 17.416 ;
			LAYER M3 ;
			RECT 60.327 17.336 60.575 17.416 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 19.352 60.575 19.432 ;
			LAYER M2 ;
			RECT 60.327 19.352 60.575 19.432 ;
			LAYER M3 ;
			RECT 60.327 19.352 60.575 19.432 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 21.368 60.575 21.448 ;
			LAYER M2 ;
			RECT 60.327 21.368 60.575 21.448 ;
			LAYER M3 ;
			RECT 60.327 21.368 60.575 21.448 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 23.384 60.575 23.464 ;
			LAYER M2 ;
			RECT 60.327 23.384 60.575 23.464 ;
			LAYER M3 ;
			RECT 60.327 23.384 60.575 23.464 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 25.400 60.575 25.480 ;
			LAYER M2 ;
			RECT 60.327 25.400 60.575 25.480 ;
			LAYER M3 ;
			RECT 60.327 25.400 60.575 25.480 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 27.416 60.575 27.496 ;
			LAYER M2 ;
			RECT 60.327 27.416 60.575 27.496 ;
			LAYER M3 ;
			RECT 60.327 27.416 60.575 27.496 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 29.432 60.575 29.512 ;
			LAYER M2 ;
			RECT 60.327 29.432 60.575 29.512 ;
			LAYER M3 ;
			RECT 60.327 29.432 60.575 29.512 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 31.448 60.575 31.528 ;
			LAYER M2 ;
			RECT 60.327 31.448 60.575 31.528 ;
			LAYER M3 ;
			RECT 60.327 31.448 60.575 31.528 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 46.328 60.575 46.408 ;
			LAYER M2 ;
			RECT 60.327 46.328 60.575 46.408 ;
			LAYER M3 ;
			RECT 60.327 46.328 60.575 46.408 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 48.344 60.575 48.424 ;
			LAYER M2 ;
			RECT 60.327 48.344 60.575 48.424 ;
			LAYER M3 ;
			RECT 60.327 48.344 60.575 48.424 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 50.360 60.575 50.440 ;
			LAYER M2 ;
			RECT 60.327 50.360 60.575 50.440 ;
			LAYER M3 ;
			RECT 60.327 50.360 60.575 50.440 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 52.376 60.575 52.456 ;
			LAYER M2 ;
			RECT 60.327 52.376 60.575 52.456 ;
			LAYER M3 ;
			RECT 60.327 52.376 60.575 52.456 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 54.392 60.575 54.472 ;
			LAYER M2 ;
			RECT 60.327 54.392 60.575 54.472 ;
			LAYER M3 ;
			RECT 60.327 54.392 60.575 54.472 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 56.408 60.575 56.488 ;
			LAYER M2 ;
			RECT 60.327 56.408 60.575 56.488 ;
			LAYER M3 ;
			RECT 60.327 56.408 60.575 56.488 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 58.424 60.575 58.504 ;
			LAYER M2 ;
			RECT 60.327 58.424 60.575 58.504 ;
			LAYER M3 ;
			RECT 60.327 58.424 60.575 58.504 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 60.440 60.575 60.520 ;
			LAYER M2 ;
			RECT 60.327 60.440 60.575 60.520 ;
			LAYER M3 ;
			RECT 60.327 60.440 60.575 60.520 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 62.456 60.575 62.536 ;
			LAYER M2 ;
			RECT 60.327 62.456 60.575 62.536 ;
			LAYER M3 ;
			RECT 60.327 62.456 60.575 62.536 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 64.472 60.575 64.552 ;
			LAYER M2 ;
			RECT 60.327 64.472 60.575 64.552 ;
			LAYER M3 ;
			RECT 60.327 64.472 60.575 64.552 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 66.488 60.575 66.568 ;
			LAYER M2 ;
			RECT 60.327 66.488 60.575 66.568 ;
			LAYER M3 ;
			RECT 60.327 66.488 60.575 66.568 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 68.504 60.575 68.584 ;
			LAYER M2 ;
			RECT 60.327 68.504 60.575 68.584 ;
			LAYER M3 ;
			RECT 60.327 68.504 60.575 68.584 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 70.520 60.575 70.600 ;
			LAYER M2 ;
			RECT 60.327 70.520 60.575 70.600 ;
			LAYER M3 ;
			RECT 60.327 70.520 60.575 70.600 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 72.536 60.575 72.616 ;
			LAYER M2 ;
			RECT 60.327 72.536 60.575 72.616 ;
			LAYER M3 ;
			RECT 60.327 72.536 60.575 72.616 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 74.552 60.575 74.632 ;
			LAYER M2 ;
			RECT 60.327 74.552 60.575 74.632 ;
			LAYER M3 ;
			RECT 60.327 74.552 60.575 74.632 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 76.568 60.575 76.648 ;
			LAYER M2 ;
			RECT 60.327 76.568 60.575 76.648 ;
			LAYER M3 ;
			RECT 60.327 76.568 60.575 76.648 ;
		END
		ANTENNADIFFAREA 0.045800 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.212400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA1 ;
		ANTENNADIFFAREA 0.045800 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.637000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.016400 LAYER VIA2 ;
		ANTENNADIFFAREA 0.045800 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.725000 LAYER M3 ;
	END Q[31]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 44.936 60.575 45.016 ;
			LAYER M2 ;
			RECT 60.327 44.936 60.575 45.016 ;
			LAYER M3 ;
			RECT 60.327 44.936 60.575 45.016 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128800 LAYER M1 ;
		ANTENNAMAXAREACAR 16.533000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.010200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.151800 LAYER M2 ;
		ANTENNAMAXAREACAR 21.415000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.263800 LAYER M3 ;
		ANTENNAMAXAREACAR 316.698000 LAYER M3 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 45.128 60.575 45.208 ;
			LAYER M2 ;
			RECT 60.327 45.128 60.575 45.208 ;
			LAYER M3 ;
			RECT 60.327 45.128 60.575 45.208 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128800 LAYER M1 ;
		ANTENNAMAXAREACAR 16.533000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.010200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.151800 LAYER M2 ;
		ANTENNAMAXAREACAR 21.415000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.012200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.263800 LAYER M3 ;
		ANTENNAMAXAREACAR 316.698000 LAYER M3 ;
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.428 60.455 1.548 ;
			LAYER M4 ;
			RECT 0.120 1.932 60.455 2.052 ;
			LAYER M4 ;
			RECT 0.120 2.184 60.455 2.304 ;
			LAYER M4 ;
			RECT 0.120 3.444 60.455 3.564 ;
			LAYER M4 ;
			RECT 0.120 3.948 60.455 4.068 ;
			LAYER M4 ;
			RECT 0.120 4.200 60.455 4.320 ;
			LAYER M4 ;
			RECT 0.120 5.460 60.455 5.580 ;
			LAYER M4 ;
			RECT 0.120 5.964 60.455 6.084 ;
			LAYER M4 ;
			RECT 0.120 6.216 60.455 6.336 ;
			LAYER M4 ;
			RECT 0.120 7.476 60.455 7.596 ;
			LAYER M4 ;
			RECT 0.120 7.980 60.455 8.100 ;
			LAYER M4 ;
			RECT 0.120 8.232 60.455 8.352 ;
			LAYER M4 ;
			RECT 0.120 9.492 60.455 9.612 ;
			LAYER M4 ;
			RECT 0.120 9.996 60.455 10.116 ;
			LAYER M4 ;
			RECT 0.120 10.248 60.455 10.368 ;
			LAYER M4 ;
			RECT 0.120 11.508 60.455 11.628 ;
			LAYER M4 ;
			RECT 0.120 12.012 60.455 12.132 ;
			LAYER M4 ;
			RECT 0.120 12.264 60.455 12.384 ;
			LAYER M4 ;
			RECT 0.120 13.524 60.455 13.644 ;
			LAYER M4 ;
			RECT 0.120 14.028 60.455 14.148 ;
			LAYER M4 ;
			RECT 0.120 14.280 60.455 14.400 ;
			LAYER M4 ;
			RECT 0.120 15.540 60.455 15.660 ;
			LAYER M4 ;
			RECT 0.120 16.044 60.455 16.164 ;
			LAYER M4 ;
			RECT 0.120 16.296 60.455 16.416 ;
			LAYER M4 ;
			RECT 0.120 17.556 60.455 17.676 ;
			LAYER M4 ;
			RECT 0.120 18.060 60.455 18.180 ;
			LAYER M4 ;
			RECT 0.120 18.312 60.455 18.432 ;
			LAYER M4 ;
			RECT 0.120 19.572 60.455 19.692 ;
			LAYER M4 ;
			RECT 0.120 20.076 60.455 20.196 ;
			LAYER M4 ;
			RECT 0.120 20.328 60.455 20.448 ;
			LAYER M4 ;
			RECT 0.120 21.588 60.455 21.708 ;
			LAYER M4 ;
			RECT 0.120 22.092 60.455 22.212 ;
			LAYER M4 ;
			RECT 0.120 22.344 60.455 22.464 ;
			LAYER M4 ;
			RECT 0.120 23.604 60.455 23.724 ;
			LAYER M4 ;
			RECT 0.120 24.108 60.455 24.228 ;
			LAYER M4 ;
			RECT 0.120 24.360 60.455 24.480 ;
			LAYER M4 ;
			RECT 0.120 25.620 60.455 25.740 ;
			LAYER M4 ;
			RECT 0.120 26.124 60.455 26.244 ;
			LAYER M4 ;
			RECT 0.120 26.376 60.455 26.496 ;
			LAYER M4 ;
			RECT 0.120 27.636 60.455 27.756 ;
			LAYER M4 ;
			RECT 0.120 28.140 60.455 28.260 ;
			LAYER M4 ;
			RECT 0.120 28.392 60.455 28.512 ;
			LAYER M4 ;
			RECT 0.120 29.652 60.455 29.772 ;
			LAYER M4 ;
			RECT 0.120 30.156 60.455 30.276 ;
			LAYER M4 ;
			RECT 0.120 30.408 60.455 30.528 ;
			LAYER M4 ;
			RECT 0.120 31.668 60.455 31.788 ;
			LAYER M4 ;
			RECT 0.120 32.172 60.455 32.292 ;
			LAYER M4 ;
			RECT 0.120 32.424 60.455 32.544 ;
			LAYER M4 ;
			RECT 0.120 33.700 60.455 33.820 ;
			LAYER M4 ;
			RECT 0.120 34.324 60.455 34.444 ;
			LAYER M4 ;
			RECT 0.120 34.730 60.455 34.850 ;
			LAYER M4 ;
			RECT 0.120 35.190 60.455 35.310 ;
			LAYER M4 ;
			RECT 0.120 35.650 60.455 35.770 ;
			LAYER M4 ;
			RECT 0.120 36.110 60.455 36.230 ;
			LAYER M4 ;
			RECT 0.120 36.340 60.455 36.460 ;
			LAYER M4 ;
			RECT 0.120 36.732 60.455 36.852 ;
			LAYER M4 ;
			RECT 0.120 37.882 60.455 38.002 ;
			LAYER M4 ;
			RECT 0.120 38.564 60.455 38.684 ;
			LAYER M4 ;
			RECT 0.120 39.476 60.455 39.596 ;
			LAYER M4 ;
			RECT 0.120 40.655 60.455 40.775 ;
			LAYER M4 ;
			RECT 0.120 41.344 60.455 41.464 ;
			LAYER M4 ;
			RECT 0.120 41.804 60.455 41.924 ;
			LAYER M4 ;
			RECT 0.120 42.680 60.455 42.800 ;
			LAYER M4 ;
			RECT 0.120 43.140 60.455 43.260 ;
			LAYER M4 ;
			RECT 0.120 44.008 60.455 44.128 ;
			LAYER M4 ;
			RECT 0.120 44.442 60.455 44.562 ;
			LAYER M4 ;
			RECT 0.120 44.902 60.455 45.022 ;
			LAYER M4 ;
			RECT 0.120 45.312 60.455 45.432 ;
			LAYER M4 ;
			RECT 0.120 45.772 60.455 45.892 ;
			LAYER M4 ;
			RECT 0.120 46.548 60.455 46.668 ;
			LAYER M4 ;
			RECT 0.120 47.052 60.455 47.172 ;
			LAYER M4 ;
			RECT 0.120 47.304 60.455 47.424 ;
			LAYER M4 ;
			RECT 0.120 48.564 60.455 48.684 ;
			LAYER M4 ;
			RECT 0.120 49.068 60.455 49.188 ;
			LAYER M4 ;
			RECT 0.120 49.320 60.455 49.440 ;
			LAYER M4 ;
			RECT 0.120 50.580 60.455 50.700 ;
			LAYER M4 ;
			RECT 0.120 51.084 60.455 51.204 ;
			LAYER M4 ;
			RECT 0.120 51.336 60.455 51.456 ;
			LAYER M4 ;
			RECT 0.120 52.596 60.455 52.716 ;
			LAYER M4 ;
			RECT 0.120 53.100 60.455 53.220 ;
			LAYER M4 ;
			RECT 0.120 53.352 60.455 53.472 ;
			LAYER M4 ;
			RECT 0.120 54.612 60.455 54.732 ;
			LAYER M4 ;
			RECT 0.120 55.116 60.455 55.236 ;
			LAYER M4 ;
			RECT 0.120 55.368 60.455 55.488 ;
			LAYER M4 ;
			RECT 0.120 56.628 60.455 56.748 ;
			LAYER M4 ;
			RECT 0.120 57.132 60.455 57.252 ;
			LAYER M4 ;
			RECT 0.120 57.384 60.455 57.504 ;
			LAYER M4 ;
			RECT 0.120 58.644 60.455 58.764 ;
			LAYER M4 ;
			RECT 0.120 59.148 60.455 59.268 ;
			LAYER M4 ;
			RECT 0.120 59.400 60.455 59.520 ;
			LAYER M4 ;
			RECT 0.120 60.660 60.455 60.780 ;
			LAYER M4 ;
			RECT 0.120 61.164 60.455 61.284 ;
			LAYER M4 ;
			RECT 0.120 61.416 60.455 61.536 ;
			LAYER M4 ;
			RECT 0.120 62.676 60.455 62.796 ;
			LAYER M4 ;
			RECT 0.120 63.180 60.455 63.300 ;
			LAYER M4 ;
			RECT 0.120 63.432 60.455 63.552 ;
			LAYER M4 ;
			RECT 0.120 64.692 60.455 64.812 ;
			LAYER M4 ;
			RECT 0.120 65.196 60.455 65.316 ;
			LAYER M4 ;
			RECT 0.120 65.448 60.455 65.568 ;
			LAYER M4 ;
			RECT 0.120 66.708 60.455 66.828 ;
			LAYER M4 ;
			RECT 0.120 67.212 60.455 67.332 ;
			LAYER M4 ;
			RECT 0.120 67.464 60.455 67.584 ;
			LAYER M4 ;
			RECT 0.120 68.724 60.455 68.844 ;
			LAYER M4 ;
			RECT 0.120 69.228 60.455 69.348 ;
			LAYER M4 ;
			RECT 0.120 69.480 60.455 69.600 ;
			LAYER M4 ;
			RECT 0.120 70.740 60.455 70.860 ;
			LAYER M4 ;
			RECT 0.120 71.244 60.455 71.364 ;
			LAYER M4 ;
			RECT 0.120 71.496 60.455 71.616 ;
			LAYER M4 ;
			RECT 0.120 72.756 60.455 72.876 ;
			LAYER M4 ;
			RECT 0.120 73.260 60.455 73.380 ;
			LAYER M4 ;
			RECT 0.120 73.512 60.455 73.632 ;
			LAYER M4 ;
			RECT 0.120 74.772 60.455 74.892 ;
			LAYER M4 ;
			RECT 0.120 75.276 60.455 75.396 ;
			LAYER M4 ;
			RECT 0.120 75.528 60.455 75.648 ;
			LAYER M4 ;
			RECT 0.120 76.788 60.455 76.908 ;
			LAYER M4 ;
			RECT 0.120 77.292 60.455 77.412 ;
			LAYER M4 ;
			RECT 0.120 77.544 60.455 77.664 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.176 60.455 1.296 ;
			LAYER M4 ;
			RECT 0.120 1.680 60.455 1.800 ;
			LAYER M4 ;
			RECT 0.120 2.688 60.455 2.808 ;
			LAYER M4 ;
			RECT 0.120 3.192 60.455 3.312 ;
			LAYER M4 ;
			RECT 0.120 3.696 60.455 3.816 ;
			LAYER M4 ;
			RECT 0.120 4.704 60.455 4.824 ;
			LAYER M4 ;
			RECT 0.120 5.208 60.455 5.328 ;
			LAYER M4 ;
			RECT 0.120 5.712 60.455 5.832 ;
			LAYER M4 ;
			RECT 0.120 6.720 60.455 6.840 ;
			LAYER M4 ;
			RECT 0.120 7.224 60.455 7.344 ;
			LAYER M4 ;
			RECT 0.120 7.728 60.455 7.848 ;
			LAYER M4 ;
			RECT 0.120 8.736 60.455 8.856 ;
			LAYER M4 ;
			RECT 0.120 9.240 60.455 9.360 ;
			LAYER M4 ;
			RECT 0.120 9.744 60.455 9.864 ;
			LAYER M4 ;
			RECT 0.120 10.752 60.455 10.872 ;
			LAYER M4 ;
			RECT 0.120 11.256 60.455 11.376 ;
			LAYER M4 ;
			RECT 0.120 11.760 60.455 11.880 ;
			LAYER M4 ;
			RECT 0.120 12.768 60.455 12.888 ;
			LAYER M4 ;
			RECT 0.120 13.272 60.455 13.392 ;
			LAYER M4 ;
			RECT 0.120 13.776 60.455 13.896 ;
			LAYER M4 ;
			RECT 0.120 14.784 60.455 14.904 ;
			LAYER M4 ;
			RECT 0.120 15.288 60.455 15.408 ;
			LAYER M4 ;
			RECT 0.120 15.792 60.455 15.912 ;
			LAYER M4 ;
			RECT 0.120 16.800 60.455 16.920 ;
			LAYER M4 ;
			RECT 0.120 17.304 60.455 17.424 ;
			LAYER M4 ;
			RECT 0.120 17.808 60.455 17.928 ;
			LAYER M4 ;
			RECT 0.120 18.816 60.455 18.936 ;
			LAYER M4 ;
			RECT 0.120 19.320 60.455 19.440 ;
			LAYER M4 ;
			RECT 0.120 19.824 60.455 19.944 ;
			LAYER M4 ;
			RECT 0.120 20.832 60.455 20.952 ;
			LAYER M4 ;
			RECT 0.120 21.336 60.455 21.456 ;
			LAYER M4 ;
			RECT 0.120 21.840 60.455 21.960 ;
			LAYER M4 ;
			RECT 0.120 22.848 60.455 22.968 ;
			LAYER M4 ;
			RECT 0.120 23.352 60.455 23.472 ;
			LAYER M4 ;
			RECT 0.120 23.856 60.455 23.976 ;
			LAYER M4 ;
			RECT 0.120 24.864 60.455 24.984 ;
			LAYER M4 ;
			RECT 0.120 25.368 60.455 25.488 ;
			LAYER M4 ;
			RECT 0.120 25.872 60.455 25.992 ;
			LAYER M4 ;
			RECT 0.120 26.880 60.455 27.000 ;
			LAYER M4 ;
			RECT 0.120 27.384 60.455 27.504 ;
			LAYER M4 ;
			RECT 0.120 27.888 60.455 28.008 ;
			LAYER M4 ;
			RECT 0.120 28.896 60.455 29.016 ;
			LAYER M4 ;
			RECT 0.120 29.400 60.455 29.520 ;
			LAYER M4 ;
			RECT 0.120 29.904 60.455 30.024 ;
			LAYER M4 ;
			RECT 0.120 30.912 60.455 31.032 ;
			LAYER M4 ;
			RECT 0.120 31.416 60.455 31.536 ;
			LAYER M4 ;
			RECT 0.120 31.920 60.455 32.040 ;
			LAYER M4 ;
			RECT 0.120 32.928 60.455 33.048 ;
			LAYER M4 ;
			RECT 0.120 34.094 60.455 34.214 ;
			LAYER M4 ;
			RECT 0.120 34.960 60.455 35.080 ;
			LAYER M4 ;
			RECT 0.120 35.420 60.455 35.540 ;
			LAYER M4 ;
			RECT 0.120 35.880 60.455 36.000 ;
			LAYER M4 ;
			RECT 0.120 36.962 60.455 37.082 ;
			LAYER M4 ;
			RECT 0.120 37.652 60.455 37.772 ;
			LAYER M4 ;
			RECT 0.120 38.794 60.455 38.914 ;
			LAYER M4 ;
			RECT 0.120 39.706 60.455 39.826 ;
			LAYER M4 ;
			RECT 0.120 40.425 60.455 40.545 ;
			LAYER M4 ;
			RECT 0.120 41.574 60.455 41.694 ;
			LAYER M4 ;
			RECT 0.120 42.034 60.455 42.154 ;
			LAYER M4 ;
			RECT 0.120 42.450 60.455 42.570 ;
			LAYER M4 ;
			RECT 0.120 42.910 60.455 43.030 ;
			LAYER M4 ;
			RECT 0.120 43.370 60.455 43.490 ;
			LAYER M4 ;
			RECT 0.120 43.778 60.455 43.898 ;
			LAYER M4 ;
			RECT 0.120 44.672 60.455 44.792 ;
			LAYER M4 ;
			RECT 0.120 45.542 60.455 45.662 ;
			LAYER M4 ;
			RECT 0.120 46.296 60.455 46.416 ;
			LAYER M4 ;
			RECT 0.120 46.800 60.455 46.920 ;
			LAYER M4 ;
			RECT 0.120 47.808 60.455 47.928 ;
			LAYER M4 ;
			RECT 0.120 48.312 60.455 48.432 ;
			LAYER M4 ;
			RECT 0.120 48.816 60.455 48.936 ;
			LAYER M4 ;
			RECT 0.120 49.824 60.455 49.944 ;
			LAYER M4 ;
			RECT 0.120 50.328 60.455 50.448 ;
			LAYER M4 ;
			RECT 0.120 50.832 60.455 50.952 ;
			LAYER M4 ;
			RECT 0.120 51.840 60.455 51.960 ;
			LAYER M4 ;
			RECT 0.120 52.344 60.455 52.464 ;
			LAYER M4 ;
			RECT 0.120 52.848 60.455 52.968 ;
			LAYER M4 ;
			RECT 0.120 53.856 60.455 53.976 ;
			LAYER M4 ;
			RECT 0.120 54.360 60.455 54.480 ;
			LAYER M4 ;
			RECT 0.120 54.864 60.455 54.984 ;
			LAYER M4 ;
			RECT 0.120 55.872 60.455 55.992 ;
			LAYER M4 ;
			RECT 0.120 56.376 60.455 56.496 ;
			LAYER M4 ;
			RECT 0.120 56.880 60.455 57.000 ;
			LAYER M4 ;
			RECT 0.120 57.888 60.455 58.008 ;
			LAYER M4 ;
			RECT 0.120 58.392 60.455 58.512 ;
			LAYER M4 ;
			RECT 0.120 58.896 60.455 59.016 ;
			LAYER M4 ;
			RECT 0.120 59.904 60.455 60.024 ;
			LAYER M4 ;
			RECT 0.120 60.408 60.455 60.528 ;
			LAYER M4 ;
			RECT 0.120 60.912 60.455 61.032 ;
			LAYER M4 ;
			RECT 0.120 61.920 60.455 62.040 ;
			LAYER M4 ;
			RECT 0.120 62.424 60.455 62.544 ;
			LAYER M4 ;
			RECT 0.120 62.928 60.455 63.048 ;
			LAYER M4 ;
			RECT 0.120 63.936 60.455 64.056 ;
			LAYER M4 ;
			RECT 0.120 64.440 60.455 64.560 ;
			LAYER M4 ;
			RECT 0.120 64.944 60.455 65.064 ;
			LAYER M4 ;
			RECT 0.120 65.952 60.455 66.072 ;
			LAYER M4 ;
			RECT 0.120 66.456 60.455 66.576 ;
			LAYER M4 ;
			RECT 0.120 66.960 60.455 67.080 ;
			LAYER M4 ;
			RECT 0.120 67.968 60.455 68.088 ;
			LAYER M4 ;
			RECT 0.120 68.472 60.455 68.592 ;
			LAYER M4 ;
			RECT 0.120 68.976 60.455 69.096 ;
			LAYER M4 ;
			RECT 0.120 69.984 60.455 70.104 ;
			LAYER M4 ;
			RECT 0.120 70.488 60.455 70.608 ;
			LAYER M4 ;
			RECT 0.120 70.992 60.455 71.112 ;
			LAYER M4 ;
			RECT 0.120 72.000 60.455 72.120 ;
			LAYER M4 ;
			RECT 0.120 72.504 60.455 72.624 ;
			LAYER M4 ;
			RECT 0.120 73.008 60.455 73.128 ;
			LAYER M4 ;
			RECT 0.120 74.016 60.455 74.136 ;
			LAYER M4 ;
			RECT 0.120 74.520 60.455 74.640 ;
			LAYER M4 ;
			RECT 0.120 75.024 60.455 75.144 ;
			LAYER M4 ;
			RECT 0.120 76.032 60.455 76.152 ;
			LAYER M4 ;
			RECT 0.120 76.536 60.455 76.656 ;
			LAYER M4 ;
			RECT 0.120 77.040 60.455 77.160 ;
			LAYER M4 ;
			RECT 0.120 78.048 60.455 78.168 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 37.832 60.575 37.912 ;
			LAYER M2 ;
			RECT 60.327 37.832 60.575 37.912 ;
			LAYER M3 ;
			RECT 60.327 37.832 60.575 37.912 ;
		END
		ANTENNAGATEAREA 0.008100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.081400 LAYER M1 ;
		ANTENNAMAXAREACAR 2.809400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.253400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.008100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.120400 LAYER M2 ;
		ANTENNAMAXAREACAR 10.990000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.507000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.008100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.163600 LAYER M3 ;
		ANTENNAMAXAREACAR 30.908400 LAYER M3 ;
	END WEB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 37.640 60.575 37.720 ;
			LAYER M2 ;
			RECT 60.327 37.640 60.575 37.720 ;
			LAYER M3 ;
			RECT 60.327 37.640 60.575 37.720 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100400 LAYER M1 ;
		ANTENNAMAXAREACAR 9.811400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.230600 LAYER M2 ;
		ANTENNAMAXAREACAR 46.438600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.855800 LAYER M3 ;
		ANTENNAMAXAREACAR 215.957000 LAYER M3 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.327 38.792 60.575 38.872 ;
			LAYER M2 ;
			RECT 60.327 38.792 60.575 38.872 ;
			LAYER M3 ;
			RECT 60.327 38.792 60.575 38.872 ;
		END
		ANTENNAGATEAREA 0.004200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.100400 LAYER M1 ;
		ANTENNAMAXAREACAR 9.811400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.483000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.004200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.230600 LAYER M2 ;
		ANTENNAMAXAREACAR 46.438600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.008200 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.966000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.004200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.855800 LAYER M3 ;
		ANTENNAMAXAREACAR 215.957000 LAYER M3 ;
	END WTSEL[1]

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 60.575 79.344 ;
		LAYER M2 ;
		RECT 0.000 0.000 60.575 79.344 ;
		LAYER M3 ;
		RECT 0.000 0.000 60.575 79.344 ;
		LAYER M4 ;
		RECT 0.276 78.793 60.175 78.913 ;
		LAYER M4 ;
		RECT 0.300 0.431 60.175 0.551 ;
		LAYER M4 ;
		RECT 0.783 45.112 58.953 45.189 ;
		LAYER M4 ;
		RECT 1.218 38.069 58.953 38.167 ;
		LAYER M4 ;
		RECT 1.218 38.249 58.953 38.347 ;
		LAYER M4 ;
		RECT 1.218 38.429 58.953 38.527 ;
		LAYER M4 ;
		RECT 1.218 38.981 58.953 39.079 ;
		LAYER M4 ;
		RECT 1.218 39.161 58.953 39.259 ;
		LAYER M4 ;
		RECT 1.218 39.341 58.953 39.439 ;
		LAYER M4 ;
		RECT 1.218 39.927 58.953 40.025 ;
		LAYER M4 ;
		RECT 1.218 40.107 58.953 40.205 ;
		LAYER M4 ;
		RECT 1.218 40.287 58.953 40.385 ;
		LAYER M4 ;
		RECT 1.218 40.839 58.953 40.937 ;
		LAYER M4 ;
		RECT 1.218 41.019 58.953 41.117 ;
		LAYER M4 ;
		RECT 1.218 41.199 58.953 41.297 ;
		LAYER M4 ;
		RECT 1.627 37.117 58.953 37.215 ;
		LAYER M4 ;
		RECT 1.627 37.297 58.953 37.395 ;
		LAYER M4 ;
		RECT 1.627 37.477 58.953 37.575 ;
		LAYER M4 ;
		RECT 51.307 1.330 52.289 1.394 ;
		LAYER M4 ;
		RECT 51.307 2.590 52.289 2.654 ;
		LAYER M4 ;
		RECT 51.307 3.346 52.289 3.410 ;
		LAYER M4 ;
		RECT 51.307 4.606 52.289 4.670 ;
		LAYER M4 ;
		RECT 51.307 5.362 52.289 5.426 ;
		LAYER M4 ;
		RECT 51.307 6.622 52.289 6.686 ;
		LAYER M4 ;
		RECT 51.307 7.378 52.289 7.442 ;
		LAYER M4 ;
		RECT 51.307 8.638 52.289 8.702 ;
		LAYER M4 ;
		RECT 51.307 9.394 52.289 9.458 ;
		LAYER M4 ;
		RECT 51.307 10.654 52.289 10.718 ;
		LAYER M4 ;
		RECT 51.307 11.410 52.289 11.474 ;
		LAYER M4 ;
		RECT 51.307 12.670 52.289 12.734 ;
		LAYER M4 ;
		RECT 51.307 13.426 52.289 13.490 ;
		LAYER M4 ;
		RECT 51.307 14.686 52.289 14.750 ;
		LAYER M4 ;
		RECT 51.307 15.442 52.289 15.506 ;
		LAYER M4 ;
		RECT 51.307 16.702 52.289 16.766 ;
		LAYER M4 ;
		RECT 51.307 17.458 52.289 17.522 ;
		LAYER M4 ;
		RECT 51.307 18.718 52.289 18.782 ;
		LAYER M4 ;
		RECT 51.307 19.474 52.289 19.538 ;
		LAYER M4 ;
		RECT 51.307 20.734 52.289 20.798 ;
		LAYER M4 ;
		RECT 51.307 21.490 52.289 21.554 ;
		LAYER M4 ;
		RECT 51.307 22.750 52.289 22.814 ;
		LAYER M4 ;
		RECT 51.307 23.506 52.289 23.570 ;
		LAYER M4 ;
		RECT 51.307 24.766 52.289 24.830 ;
		LAYER M4 ;
		RECT 51.307 25.522 52.289 25.586 ;
		LAYER M4 ;
		RECT 51.307 26.782 52.289 26.846 ;
		LAYER M4 ;
		RECT 51.307 27.538 52.289 27.602 ;
		LAYER M4 ;
		RECT 51.307 28.798 52.289 28.862 ;
		LAYER M4 ;
		RECT 51.307 29.554 52.289 29.618 ;
		LAYER M4 ;
		RECT 51.307 30.814 52.289 30.878 ;
		LAYER M4 ;
		RECT 51.307 31.570 52.289 31.634 ;
		LAYER M4 ;
		RECT 51.307 32.830 52.289 32.894 ;
		LAYER M4 ;
		RECT 51.307 46.450 52.289 46.514 ;
		LAYER M4 ;
		RECT 51.307 47.710 52.289 47.774 ;
		LAYER M4 ;
		RECT 51.307 48.466 52.289 48.530 ;
		LAYER M4 ;
		RECT 51.307 49.726 52.289 49.790 ;
		LAYER M4 ;
		RECT 51.307 50.482 52.289 50.546 ;
		LAYER M4 ;
		RECT 51.307 51.742 52.289 51.806 ;
		LAYER M4 ;
		RECT 51.307 52.498 52.289 52.562 ;
		LAYER M4 ;
		RECT 51.307 53.758 52.289 53.822 ;
		LAYER M4 ;
		RECT 51.307 54.514 52.289 54.578 ;
		LAYER M4 ;
		RECT 51.307 55.774 52.289 55.838 ;
		LAYER M4 ;
		RECT 51.307 56.530 52.289 56.594 ;
		LAYER M4 ;
		RECT 51.307 57.790 52.289 57.854 ;
		LAYER M4 ;
		RECT 51.307 58.546 52.289 58.610 ;
		LAYER M4 ;
		RECT 51.307 59.806 52.289 59.870 ;
		LAYER M4 ;
		RECT 51.307 60.562 52.289 60.626 ;
		LAYER M4 ;
		RECT 51.307 61.822 52.289 61.886 ;
		LAYER M4 ;
		RECT 51.307 62.578 52.289 62.642 ;
		LAYER M4 ;
		RECT 51.307 63.838 52.289 63.902 ;
		LAYER M4 ;
		RECT 51.307 64.594 52.289 64.658 ;
		LAYER M4 ;
		RECT 51.307 65.854 52.289 65.918 ;
		LAYER M4 ;
		RECT 51.307 66.610 52.289 66.674 ;
		LAYER M4 ;
		RECT 51.307 67.870 52.289 67.934 ;
		LAYER M4 ;
		RECT 51.307 68.626 52.289 68.690 ;
		LAYER M4 ;
		RECT 51.307 69.886 52.289 69.950 ;
		LAYER M4 ;
		RECT 51.307 70.642 52.289 70.706 ;
		LAYER M4 ;
		RECT 51.307 71.902 52.289 71.966 ;
		LAYER M4 ;
		RECT 51.307 72.658 52.289 72.722 ;
		LAYER M4 ;
		RECT 51.307 73.918 52.289 73.982 ;
		LAYER M4 ;
		RECT 51.307 74.674 52.289 74.738 ;
		LAYER M4 ;
		RECT 51.307 75.934 52.289 75.998 ;
		LAYER M4 ;
		RECT 51.307 76.690 52.289 76.754 ;
		LAYER M4 ;
		RECT 51.307 77.950 52.289 78.014 ;
		LAYER M4 ;
		RECT 52.816 1.337 54.539 1.387 ;
		LAYER M4 ;
		RECT 52.816 2.597 54.731 2.647 ;
		LAYER M4 ;
		RECT 52.816 3.353 54.539 3.403 ;
		LAYER M4 ;
		RECT 52.816 4.613 54.731 4.663 ;
		LAYER M4 ;
		RECT 52.816 5.369 54.539 5.419 ;
		LAYER M4 ;
		RECT 52.816 6.629 54.731 6.679 ;
		LAYER M4 ;
		RECT 52.816 7.385 54.539 7.435 ;
		LAYER M4 ;
		RECT 52.816 8.645 54.731 8.695 ;
		LAYER M4 ;
		RECT 52.816 9.401 54.539 9.451 ;
		LAYER M4 ;
		RECT 52.816 10.661 54.731 10.711 ;
		LAYER M4 ;
		RECT 52.816 11.417 54.539 11.467 ;
		LAYER M4 ;
		RECT 52.816 12.677 54.731 12.727 ;
		LAYER M4 ;
		RECT 52.816 13.433 54.539 13.483 ;
		LAYER M4 ;
		RECT 52.816 14.693 54.731 14.743 ;
		LAYER M4 ;
		RECT 52.816 15.449 54.539 15.499 ;
		LAYER M4 ;
		RECT 52.816 16.709 54.731 16.759 ;
		LAYER M4 ;
		RECT 52.816 17.465 54.539 17.515 ;
		LAYER M4 ;
		RECT 52.816 18.725 54.731 18.775 ;
		LAYER M4 ;
		RECT 52.816 19.481 54.539 19.531 ;
		LAYER M4 ;
		RECT 52.816 20.741 54.731 20.791 ;
		LAYER M4 ;
		RECT 52.816 21.497 54.539 21.547 ;
		LAYER M4 ;
		RECT 52.816 22.757 54.731 22.807 ;
		LAYER M4 ;
		RECT 52.816 23.513 54.539 23.563 ;
		LAYER M4 ;
		RECT 52.816 24.773 54.731 24.823 ;
		LAYER M4 ;
		RECT 52.816 25.529 54.539 25.579 ;
		LAYER M4 ;
		RECT 52.816 26.789 54.731 26.839 ;
		LAYER M4 ;
		RECT 52.816 27.545 54.539 27.595 ;
		LAYER M4 ;
		RECT 52.816 28.805 54.731 28.855 ;
		LAYER M4 ;
		RECT 52.816 29.561 54.539 29.611 ;
		LAYER M4 ;
		RECT 52.816 30.821 54.731 30.871 ;
		LAYER M4 ;
		RECT 52.816 31.577 54.539 31.627 ;
		LAYER M4 ;
		RECT 52.816 32.837 54.731 32.887 ;
		LAYER M4 ;
		RECT 52.816 46.457 54.539 46.507 ;
		LAYER M4 ;
		RECT 52.816 47.717 54.731 47.767 ;
		LAYER M4 ;
		RECT 52.816 48.473 54.539 48.523 ;
		LAYER M4 ;
		RECT 52.816 49.733 54.731 49.783 ;
		LAYER M4 ;
		RECT 52.816 50.489 54.539 50.539 ;
		LAYER M4 ;
		RECT 52.816 51.749 54.731 51.799 ;
		LAYER M4 ;
		RECT 52.816 52.505 54.539 52.555 ;
		LAYER M4 ;
		RECT 52.816 53.765 54.731 53.815 ;
		LAYER M4 ;
		RECT 52.816 54.521 54.539 54.571 ;
		LAYER M4 ;
		RECT 52.816 55.781 54.731 55.831 ;
		LAYER M4 ;
		RECT 52.816 56.537 54.539 56.587 ;
		LAYER M4 ;
		RECT 52.816 57.797 54.731 57.847 ;
		LAYER M4 ;
		RECT 52.816 58.553 54.539 58.603 ;
		LAYER M4 ;
		RECT 52.816 59.813 54.731 59.863 ;
		LAYER M4 ;
		RECT 52.816 60.569 54.539 60.619 ;
		LAYER M4 ;
		RECT 52.816 61.829 54.731 61.879 ;
		LAYER M4 ;
		RECT 52.816 62.585 54.539 62.635 ;
		LAYER M4 ;
		RECT 52.816 63.845 54.731 63.895 ;
		LAYER M4 ;
		RECT 52.816 64.601 54.539 64.651 ;
		LAYER M4 ;
		RECT 52.816 65.861 54.731 65.911 ;
		LAYER M4 ;
		RECT 52.816 66.617 54.539 66.667 ;
		LAYER M4 ;
		RECT 52.816 67.877 54.731 67.927 ;
		LAYER M4 ;
		RECT 52.816 68.633 54.539 68.683 ;
		LAYER M4 ;
		RECT 52.816 69.893 54.731 69.943 ;
		LAYER M4 ;
		RECT 52.816 70.649 54.539 70.699 ;
		LAYER M4 ;
		RECT 52.816 71.909 54.731 71.959 ;
		LAYER M4 ;
		RECT 52.816 72.665 54.539 72.715 ;
		LAYER M4 ;
		RECT 52.816 73.925 54.731 73.975 ;
		LAYER M4 ;
		RECT 52.816 74.681 54.539 74.731 ;
		LAYER M4 ;
		RECT 52.816 75.941 54.731 75.991 ;
		LAYER M4 ;
		RECT 52.816 76.697 54.539 76.747 ;
		LAYER M4 ;
		RECT 52.816 77.957 54.731 78.007 ;
		LAYER M4 ;
		RECT 53.917 1.589 54.809 1.639 ;
		LAYER M4 ;
		RECT 53.917 2.345 54.809 2.395 ;
		LAYER M4 ;
		RECT 53.917 3.605 54.809 3.655 ;
		LAYER M4 ;
		RECT 53.917 4.361 54.809 4.411 ;
		LAYER M4 ;
		RECT 53.917 5.621 54.809 5.671 ;
		LAYER M4 ;
		RECT 53.917 6.377 54.809 6.427 ;
		LAYER M4 ;
		RECT 53.917 7.637 54.809 7.687 ;
		LAYER M4 ;
		RECT 53.917 8.393 54.809 8.443 ;
		LAYER M4 ;
		RECT 53.917 9.653 54.809 9.703 ;
		LAYER M4 ;
		RECT 53.917 10.409 54.809 10.459 ;
		LAYER M4 ;
		RECT 53.917 11.669 54.809 11.719 ;
		LAYER M4 ;
		RECT 53.917 12.425 54.809 12.475 ;
		LAYER M4 ;
		RECT 53.917 13.685 54.809 13.735 ;
		LAYER M4 ;
		RECT 53.917 14.441 54.809 14.491 ;
		LAYER M4 ;
		RECT 53.917 15.701 54.809 15.751 ;
		LAYER M4 ;
		RECT 53.917 16.457 54.809 16.507 ;
		LAYER M4 ;
		RECT 53.917 17.717 54.809 17.767 ;
		LAYER M4 ;
		RECT 53.917 18.473 54.809 18.523 ;
		LAYER M4 ;
		RECT 53.917 19.733 54.809 19.783 ;
		LAYER M4 ;
		RECT 53.917 20.489 54.809 20.539 ;
		LAYER M4 ;
		RECT 53.917 21.749 54.809 21.799 ;
		LAYER M4 ;
		RECT 53.917 22.505 54.809 22.555 ;
		LAYER M4 ;
		RECT 53.917 23.765 54.809 23.815 ;
		LAYER M4 ;
		RECT 53.917 24.521 54.809 24.571 ;
		LAYER M4 ;
		RECT 53.917 25.781 54.809 25.831 ;
		LAYER M4 ;
		RECT 53.917 26.537 54.809 26.587 ;
		LAYER M4 ;
		RECT 53.917 27.797 54.809 27.847 ;
		LAYER M4 ;
		RECT 53.917 28.553 54.809 28.603 ;
		LAYER M4 ;
		RECT 53.917 29.813 54.809 29.863 ;
		LAYER M4 ;
		RECT 53.917 30.569 54.809 30.619 ;
		LAYER M4 ;
		RECT 53.917 31.829 54.809 31.879 ;
		LAYER M4 ;
		RECT 53.917 32.585 54.809 32.635 ;
		LAYER M4 ;
		RECT 53.917 46.709 54.809 46.759 ;
		LAYER M4 ;
		RECT 53.917 47.465 54.809 47.515 ;
		LAYER M4 ;
		RECT 53.917 48.725 54.809 48.775 ;
		LAYER M4 ;
		RECT 53.917 49.481 54.809 49.531 ;
		LAYER M4 ;
		RECT 53.917 50.741 54.809 50.791 ;
		LAYER M4 ;
		RECT 53.917 51.497 54.809 51.547 ;
		LAYER M4 ;
		RECT 53.917 52.757 54.809 52.807 ;
		LAYER M4 ;
		RECT 53.917 53.513 54.809 53.563 ;
		LAYER M4 ;
		RECT 53.917 54.773 54.809 54.823 ;
		LAYER M4 ;
		RECT 53.917 55.529 54.809 55.579 ;
		LAYER M4 ;
		RECT 53.917 56.789 54.809 56.839 ;
		LAYER M4 ;
		RECT 53.917 57.545 54.809 57.595 ;
		LAYER M4 ;
		RECT 53.917 58.805 54.809 58.855 ;
		LAYER M4 ;
		RECT 53.917 59.561 54.809 59.611 ;
		LAYER M4 ;
		RECT 53.917 60.821 54.809 60.871 ;
		LAYER M4 ;
		RECT 53.917 61.577 54.809 61.627 ;
		LAYER M4 ;
		RECT 53.917 62.837 54.809 62.887 ;
		LAYER M4 ;
		RECT 53.917 63.593 54.809 63.643 ;
		LAYER M4 ;
		RECT 53.917 64.853 54.809 64.903 ;
		LAYER M4 ;
		RECT 53.917 65.609 54.809 65.659 ;
		LAYER M4 ;
		RECT 53.917 66.869 54.809 66.919 ;
		LAYER M4 ;
		RECT 53.917 67.625 54.809 67.675 ;
		LAYER M4 ;
		RECT 53.917 68.885 54.809 68.935 ;
		LAYER M4 ;
		RECT 53.917 69.641 54.809 69.691 ;
		LAYER M4 ;
		RECT 53.917 70.901 54.809 70.951 ;
		LAYER M4 ;
		RECT 53.917 71.657 54.809 71.707 ;
		LAYER M4 ;
		RECT 53.917 72.917 54.809 72.967 ;
		LAYER M4 ;
		RECT 53.917 73.673 54.809 73.723 ;
		LAYER M4 ;
		RECT 53.917 74.933 54.809 74.983 ;
		LAYER M4 ;
		RECT 53.917 75.689 54.809 75.739 ;
		LAYER M4 ;
		RECT 53.917 76.949 54.809 76.999 ;
		LAYER M4 ;
		RECT 53.917 77.705 54.809 77.755 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 60.575 79.344 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 60.575 79.344 ;
	END
END TS1N16FFCLLSVTA1024X32M4SW

END LIBRARY
