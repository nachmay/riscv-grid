# Created by MC2 : Version 2013.12.00.f on 2025/06/23, 08:27:50

#*********************************************************************************************************************/
# Technology     : TSMC 16nm CMOS Logic FinFet Compact (FFC) Low Leakage HKMG                          */
# Memory Type    : TSMC 16nm FFC Single Port SRAM with d0907 bit cell                     */
# Library Name   : ts1n16ffcllsvta8192x32m8sw (user specify : ts1n16ffcllsvta8192x32m8sw)            */
# Library Version: 120a                                                */
# Generated Time : 2025/06/23, 08:27:44                                        */
#*********************************************************************************************************************/
#                                                            */
# STATEMENT OF USE                                                    */
#                                                            */
# This information contains confidential and proprietary information of TSMC.                    */
# No part of this information may be reproduced, transmitted, transcribed,                        */
# stored in a retrieval system, or translated into any human or computer                        */
# language, in any form or by any means, electronic, mechanical, magnetic,                        */
# optical, chemical, manual, or otherwise, without the prior written permission                    */
# of TSMC. This information was prepared for informational purpose and is for                    */
# use by TSMC's customers only. TSMC reserves the right to make changes in the                    */
# information at any time and without notice.                                    */
#                                                            */
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N16FFCLLSVTA8192X32M8SW
	CLASS BLOCK ;
	FOREIGN TS1N16FFCLLSVTA8192X32M8SW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 220.677 BY 144.672 ;
	SYMMETRY X Y ;
	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 63.794 220.677 63.892 ;
			LAYER M2 ;
			RECT 220.477 63.794 220.677 63.892 ;
			LAYER M3 ;
			RECT 220.477 63.794 220.677 63.892 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 64.766 220.677 64.864 ;
			LAYER M2 ;
			RECT 220.477 64.766 220.677 64.864 ;
			LAYER M3 ;
			RECT 220.477 64.766 220.677 64.864 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 66.891 220.677 66.989 ;
			LAYER M2 ;
			RECT 220.477 66.891 220.677 66.989 ;
			LAYER M3 ;
			RECT 220.477 66.891 220.677 66.989 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 69.513 220.677 69.611 ;
			LAYER M2 ;
			RECT 220.477 69.513 220.677 69.611 ;
			LAYER M3 ;
			RECT 220.477 69.513 220.677 69.611 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 69.979 220.677 70.077 ;
			LAYER M2 ;
			RECT 220.477 69.979 220.677 70.077 ;
			LAYER M3 ;
			RECT 220.477 69.979 220.677 70.077 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 76.743 220.677 76.841 ;
			LAYER M2 ;
			RECT 220.477 76.743 220.677 76.841 ;
			LAYER M3 ;
			RECT 220.477 76.743 220.677 76.841 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 70.973 220.677 71.071 ;
			LAYER M2 ;
			RECT 220.477 70.973 220.677 71.071 ;
			LAYER M3 ;
			RECT 220.477 70.973 220.677 71.071 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 71.955 220.677 72.053 ;
			LAYER M2 ;
			RECT 220.477 71.955 220.677 72.053 ;
			LAYER M3 ;
			RECT 220.477 71.955 220.677 72.053 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 72.661 220.677 72.759 ;
			LAYER M2 ;
			RECT 220.477 72.661 220.677 72.759 ;
			LAYER M3 ;
			RECT 220.477 72.661 220.677 72.759 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 74.369 220.677 74.467 ;
			LAYER M2 ;
			RECT 220.477 74.369 220.677 74.467 ;
			LAYER M3 ;
			RECT 220.477 74.369 220.677 74.467 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[9]

	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 75.147 220.677 75.245 ;
			LAYER M2 ;
			RECT 220.477 75.147 220.677 75.245 ;
			LAYER M3 ;
			RECT 220.477 75.147 220.677 75.245 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[10]

	PIN A[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 76.267 220.677 76.365 ;
			LAYER M2 ;
			RECT 220.477 76.267 220.677 76.365 ;
			LAYER M3 ;
			RECT 220.477 76.267 220.677 76.365 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[11]

	PIN A[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 78.053 220.677 78.151 ;
			LAYER M2 ;
			RECT 220.477 78.053 220.677 78.151 ;
			LAYER M3 ;
			RECT 220.477 78.053 220.677 78.151 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.163800 LAYER M1 ;
		ANTENNAMAXAREACAR 15.340900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088320 LAYER M2 ;
		ANTENNAMAXAREACAR 24.311600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.598440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.151200 LAYER M3 ;
		ANTENNAMAXAREACAR 36.752800 LAYER M3 ;
	END A[12]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 3.647 220.677 3.745 ;
			LAYER M2 ;
			RECT 220.477 3.647 220.677 3.745 ;
			LAYER M3 ;
			RECT 220.477 3.647 220.677 3.745 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 7.679 220.677 7.777 ;
			LAYER M2 ;
			RECT 220.477 7.679 220.677 7.777 ;
			LAYER M3 ;
			RECT 220.477 7.679 220.677 7.777 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 11.711 220.677 11.809 ;
			LAYER M2 ;
			RECT 220.477 11.711 220.677 11.809 ;
			LAYER M3 ;
			RECT 220.477 11.711 220.677 11.809 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 15.743 220.677 15.841 ;
			LAYER M2 ;
			RECT 220.477 15.743 220.677 15.841 ;
			LAYER M3 ;
			RECT 220.477 15.743 220.677 15.841 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 19.775 220.677 19.873 ;
			LAYER M2 ;
			RECT 220.477 19.775 220.677 19.873 ;
			LAYER M3 ;
			RECT 220.477 19.775 220.677 19.873 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 23.807 220.677 23.905 ;
			LAYER M2 ;
			RECT 220.477 23.807 220.677 23.905 ;
			LAYER M3 ;
			RECT 220.477 23.807 220.677 23.905 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 27.839 220.677 27.937 ;
			LAYER M2 ;
			RECT 220.477 27.839 220.677 27.937 ;
			LAYER M3 ;
			RECT 220.477 27.839 220.677 27.937 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 31.871 220.677 31.969 ;
			LAYER M2 ;
			RECT 220.477 31.871 220.677 31.969 ;
			LAYER M3 ;
			RECT 220.477 31.871 220.677 31.969 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 35.903 220.677 36.001 ;
			LAYER M2 ;
			RECT 220.477 35.903 220.677 36.001 ;
			LAYER M3 ;
			RECT 220.477 35.903 220.677 36.001 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 39.935 220.677 40.033 ;
			LAYER M2 ;
			RECT 220.477 39.935 220.677 40.033 ;
			LAYER M3 ;
			RECT 220.477 39.935 220.677 40.033 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 43.967 220.677 44.065 ;
			LAYER M2 ;
			RECT 220.477 43.967 220.677 44.065 ;
			LAYER M3 ;
			RECT 220.477 43.967 220.677 44.065 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 47.999 220.677 48.097 ;
			LAYER M2 ;
			RECT 220.477 47.999 220.677 48.097 ;
			LAYER M3 ;
			RECT 220.477 47.999 220.677 48.097 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 52.031 220.677 52.129 ;
			LAYER M2 ;
			RECT 220.477 52.031 220.677 52.129 ;
			LAYER M3 ;
			RECT 220.477 52.031 220.677 52.129 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 56.063 220.677 56.161 ;
			LAYER M2 ;
			RECT 220.477 56.063 220.677 56.161 ;
			LAYER M3 ;
			RECT 220.477 56.063 220.677 56.161 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 59.087 220.677 59.185 ;
			LAYER M2 ;
			RECT 220.477 59.087 220.677 59.185 ;
			LAYER M3 ;
			RECT 220.477 59.087 220.677 59.185 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 61.103 220.677 61.201 ;
			LAYER M2 ;
			RECT 220.477 61.103 220.677 61.201 ;
			LAYER M3 ;
			RECT 220.477 61.103 220.677 61.201 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 84.807 220.677 84.905 ;
			LAYER M2 ;
			RECT 220.477 84.807 220.677 84.905 ;
			LAYER M3 ;
			RECT 220.477 84.807 220.677 84.905 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 86.927 220.677 87.025 ;
			LAYER M2 ;
			RECT 220.477 86.927 220.677 87.025 ;
			LAYER M3 ;
			RECT 220.477 86.927 220.677 87.025 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 89.951 220.677 90.049 ;
			LAYER M2 ;
			RECT 220.477 89.951 220.677 90.049 ;
			LAYER M3 ;
			RECT 220.477 89.951 220.677 90.049 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 93.983 220.677 94.081 ;
			LAYER M2 ;
			RECT 220.477 93.983 220.677 94.081 ;
			LAYER M3 ;
			RECT 220.477 93.983 220.677 94.081 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 98.015 220.677 98.113 ;
			LAYER M2 ;
			RECT 220.477 98.015 220.677 98.113 ;
			LAYER M3 ;
			RECT 220.477 98.015 220.677 98.113 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 102.047 220.677 102.145 ;
			LAYER M2 ;
			RECT 220.477 102.047 220.677 102.145 ;
			LAYER M3 ;
			RECT 220.477 102.047 220.677 102.145 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 106.079 220.677 106.177 ;
			LAYER M2 ;
			RECT 220.477 106.079 220.677 106.177 ;
			LAYER M3 ;
			RECT 220.477 106.079 220.677 106.177 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 110.111 220.677 110.209 ;
			LAYER M2 ;
			RECT 220.477 110.111 220.677 110.209 ;
			LAYER M3 ;
			RECT 220.477 110.111 220.677 110.209 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 114.143 220.677 114.241 ;
			LAYER M2 ;
			RECT 220.477 114.143 220.677 114.241 ;
			LAYER M3 ;
			RECT 220.477 114.143 220.677 114.241 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 118.175 220.677 118.273 ;
			LAYER M2 ;
			RECT 220.477 118.175 220.677 118.273 ;
			LAYER M3 ;
			RECT 220.477 118.175 220.677 118.273 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 122.207 220.677 122.305 ;
			LAYER M2 ;
			RECT 220.477 122.207 220.677 122.305 ;
			LAYER M3 ;
			RECT 220.477 122.207 220.677 122.305 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 126.239 220.677 126.337 ;
			LAYER M2 ;
			RECT 220.477 126.239 220.677 126.337 ;
			LAYER M3 ;
			RECT 220.477 126.239 220.677 126.337 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 130.271 220.677 130.369 ;
			LAYER M2 ;
			RECT 220.477 130.271 220.677 130.369 ;
			LAYER M3 ;
			RECT 220.477 130.271 220.677 130.369 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 134.303 220.677 134.401 ;
			LAYER M2 ;
			RECT 220.477 134.303 220.677 134.401 ;
			LAYER M3 ;
			RECT 220.477 134.303 220.677 134.401 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 138.335 220.677 138.433 ;
			LAYER M2 ;
			RECT 220.477 138.335 220.677 138.433 ;
			LAYER M3 ;
			RECT 220.477 138.335 220.677 138.433 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 142.367 220.677 142.465 ;
			LAYER M2 ;
			RECT 220.477 142.367 220.677 142.465 ;
			LAYER M3 ;
			RECT 220.477 142.367 220.677 142.465 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.119280 LAYER M1 ;
		ANTENNAMAXAREACAR 36.498600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.106440 LAYER M2 ;
		ANTENNAMAXAREACAR 43.429700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.118920 LAYER M3 ;
		ANTENNAMAXAREACAR 74.700000 LAYER M3 ;
	END BWEB[31]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 65.787 220.677 65.885 ;
			LAYER M2 ;
			RECT 220.477 65.787 220.677 65.885 ;
			LAYER M3 ;
			RECT 220.477 65.787 220.677 65.885 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.130320 LAYER M1 ;
		ANTENNAMAXAREACAR 9.525960 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.049080 LAYER M2 ;
		ANTENNAMAXAREACAR 11.142800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.399000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.119760 LAYER M3 ;
		ANTENNAMAXAREACAR 30.577400 LAYER M3 ;
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 77.219 220.677 77.317 ;
			LAYER M2 ;
			RECT 220.477 77.219 220.677 77.317 ;
			LAYER M3 ;
			RECT 220.477 77.219 220.677 77.317 ;
		END
		ANTENNAGATEAREA 0.187200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 1.224720 LAYER M1 ;
		ANTENNAMAXAREACAR 15.343400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.040560 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.187200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 2.779200 LAYER M2 ;
		ANTENNAMAXAREACAR 431.180000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.014760 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.588920 LAYER VIA2 ;
		ANTENNAGATEAREA 0.187200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 2.196960 LAYER M3 ;
		ANTENNAMAXAREACAR 440.815000 LAYER M3 ;
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 2.313 220.677 2.411 ;
			LAYER M2 ;
			RECT 220.477 2.313 220.677 2.411 ;
			LAYER M3 ;
			RECT 220.477 2.313 220.677 2.411 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 6.345 220.677 6.443 ;
			LAYER M2 ;
			RECT 220.477 6.345 220.677 6.443 ;
			LAYER M3 ;
			RECT 220.477 6.345 220.677 6.443 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 10.377 220.677 10.475 ;
			LAYER M2 ;
			RECT 220.477 10.377 220.677 10.475 ;
			LAYER M3 ;
			RECT 220.477 10.377 220.677 10.475 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 14.409 220.677 14.507 ;
			LAYER M2 ;
			RECT 220.477 14.409 220.677 14.507 ;
			LAYER M3 ;
			RECT 220.477 14.409 220.677 14.507 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 18.441 220.677 18.539 ;
			LAYER M2 ;
			RECT 220.477 18.441 220.677 18.539 ;
			LAYER M3 ;
			RECT 220.477 18.441 220.677 18.539 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 22.473 220.677 22.571 ;
			LAYER M2 ;
			RECT 220.477 22.473 220.677 22.571 ;
			LAYER M3 ;
			RECT 220.477 22.473 220.677 22.571 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 26.505 220.677 26.603 ;
			LAYER M2 ;
			RECT 220.477 26.505 220.677 26.603 ;
			LAYER M3 ;
			RECT 220.477 26.505 220.677 26.603 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 30.537 220.677 30.635 ;
			LAYER M2 ;
			RECT 220.477 30.537 220.677 30.635 ;
			LAYER M3 ;
			RECT 220.477 30.537 220.677 30.635 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 34.569 220.677 34.667 ;
			LAYER M2 ;
			RECT 220.477 34.569 220.677 34.667 ;
			LAYER M3 ;
			RECT 220.477 34.569 220.677 34.667 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 38.601 220.677 38.699 ;
			LAYER M2 ;
			RECT 220.477 38.601 220.677 38.699 ;
			LAYER M3 ;
			RECT 220.477 38.601 220.677 38.699 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 42.633 220.677 42.731 ;
			LAYER M2 ;
			RECT 220.477 42.633 220.677 42.731 ;
			LAYER M3 ;
			RECT 220.477 42.633 220.677 42.731 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 46.665 220.677 46.763 ;
			LAYER M2 ;
			RECT 220.477 46.665 220.677 46.763 ;
			LAYER M3 ;
			RECT 220.477 46.665 220.677 46.763 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 50.697 220.677 50.795 ;
			LAYER M2 ;
			RECT 220.477 50.697 220.677 50.795 ;
			LAYER M3 ;
			RECT 220.477 50.697 220.677 50.795 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 54.729 220.677 54.827 ;
			LAYER M2 ;
			RECT 220.477 54.729 220.677 54.827 ;
			LAYER M3 ;
			RECT 220.477 54.729 220.677 54.827 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 57.753 220.677 57.851 ;
			LAYER M2 ;
			RECT 220.477 57.753 220.677 57.851 ;
			LAYER M3 ;
			RECT 220.477 57.753 220.677 57.851 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 59.769 220.677 59.867 ;
			LAYER M2 ;
			RECT 220.477 59.769 220.677 59.867 ;
			LAYER M3 ;
			RECT 220.477 59.769 220.677 59.867 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 83.537 220.677 83.635 ;
			LAYER M2 ;
			RECT 220.477 83.537 220.677 83.635 ;
			LAYER M3 ;
			RECT 220.477 83.537 220.677 83.635 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 85.593 220.677 85.691 ;
			LAYER M2 ;
			RECT 220.477 85.593 220.677 85.691 ;
			LAYER M3 ;
			RECT 220.477 85.593 220.677 85.691 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 88.617 220.677 88.715 ;
			LAYER M2 ;
			RECT 220.477 88.617 220.677 88.715 ;
			LAYER M3 ;
			RECT 220.477 88.617 220.677 88.715 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 92.649 220.677 92.747 ;
			LAYER M2 ;
			RECT 220.477 92.649 220.677 92.747 ;
			LAYER M3 ;
			RECT 220.477 92.649 220.677 92.747 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 96.681 220.677 96.779 ;
			LAYER M2 ;
			RECT 220.477 96.681 220.677 96.779 ;
			LAYER M3 ;
			RECT 220.477 96.681 220.677 96.779 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 100.713 220.677 100.811 ;
			LAYER M2 ;
			RECT 220.477 100.713 220.677 100.811 ;
			LAYER M3 ;
			RECT 220.477 100.713 220.677 100.811 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 104.745 220.677 104.843 ;
			LAYER M2 ;
			RECT 220.477 104.745 220.677 104.843 ;
			LAYER M3 ;
			RECT 220.477 104.745 220.677 104.843 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 108.777 220.677 108.875 ;
			LAYER M2 ;
			RECT 220.477 108.777 220.677 108.875 ;
			LAYER M3 ;
			RECT 220.477 108.777 220.677 108.875 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 112.809 220.677 112.907 ;
			LAYER M2 ;
			RECT 220.477 112.809 220.677 112.907 ;
			LAYER M3 ;
			RECT 220.477 112.809 220.677 112.907 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 116.841 220.677 116.939 ;
			LAYER M2 ;
			RECT 220.477 116.841 220.677 116.939 ;
			LAYER M3 ;
			RECT 220.477 116.841 220.677 116.939 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 120.873 220.677 120.971 ;
			LAYER M2 ;
			RECT 220.477 120.873 220.677 120.971 ;
			LAYER M3 ;
			RECT 220.477 120.873 220.677 120.971 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 124.905 220.677 125.003 ;
			LAYER M2 ;
			RECT 220.477 124.905 220.677 125.003 ;
			LAYER M3 ;
			RECT 220.477 124.905 220.677 125.003 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 128.937 220.677 129.035 ;
			LAYER M2 ;
			RECT 220.477 128.937 220.677 129.035 ;
			LAYER M3 ;
			RECT 220.477 128.937 220.677 129.035 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 132.969 220.677 133.067 ;
			LAYER M2 ;
			RECT 220.477 132.969 220.677 133.067 ;
			LAYER M3 ;
			RECT 220.477 132.969 220.677 133.067 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 137.001 220.677 137.099 ;
			LAYER M2 ;
			RECT 220.477 137.001 220.677 137.099 ;
			LAYER M3 ;
			RECT 220.477 137.001 220.677 137.099 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 141.033 220.677 141.131 ;
			LAYER M2 ;
			RECT 220.477 141.033 220.677 141.131 ;
			LAYER M3 ;
			RECT 220.477 141.033 220.677 141.131 ;
		END
		ANTENNAGATEAREA 0.002300 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.124080 LAYER M1 ;
		ANTENNAMAXAREACAR 34.024100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.529680 LAYER VIA1 ;
		ANTENNAGATEAREA 0.002300 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.057720 LAYER M2 ;
		ANTENNAMAXAREACAR 38.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.003720 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA2 ;
		ANTENNAGATEAREA 0.002300 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.094200 LAYER M3 ;
		ANTENNAMAXAREACAR 65.998900 LAYER M3 ;
	END D[31]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 2.075 220.677 2.173 ;
			LAYER M2 ;
			RECT 220.477 2.075 220.677 2.173 ;
			LAYER M3 ;
			RECT 220.477 2.075 220.677 2.173 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 6.107 220.677 6.205 ;
			LAYER M2 ;
			RECT 220.477 6.107 220.677 6.205 ;
			LAYER M3 ;
			RECT 220.477 6.107 220.677 6.205 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 10.139 220.677 10.237 ;
			LAYER M2 ;
			RECT 220.477 10.139 220.677 10.237 ;
			LAYER M3 ;
			RECT 220.477 10.139 220.677 10.237 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 14.171 220.677 14.269 ;
			LAYER M2 ;
			RECT 220.477 14.171 220.677 14.269 ;
			LAYER M3 ;
			RECT 220.477 14.171 220.677 14.269 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 18.203 220.677 18.301 ;
			LAYER M2 ;
			RECT 220.477 18.203 220.677 18.301 ;
			LAYER M3 ;
			RECT 220.477 18.203 220.677 18.301 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 22.235 220.677 22.333 ;
			LAYER M2 ;
			RECT 220.477 22.235 220.677 22.333 ;
			LAYER M3 ;
			RECT 220.477 22.235 220.677 22.333 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 26.267 220.677 26.365 ;
			LAYER M2 ;
			RECT 220.477 26.267 220.677 26.365 ;
			LAYER M3 ;
			RECT 220.477 26.267 220.677 26.365 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 30.299 220.677 30.397 ;
			LAYER M2 ;
			RECT 220.477 30.299 220.677 30.397 ;
			LAYER M3 ;
			RECT 220.477 30.299 220.677 30.397 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 34.331 220.677 34.429 ;
			LAYER M2 ;
			RECT 220.477 34.331 220.677 34.429 ;
			LAYER M3 ;
			RECT 220.477 34.331 220.677 34.429 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 38.363 220.677 38.461 ;
			LAYER M2 ;
			RECT 220.477 38.363 220.677 38.461 ;
			LAYER M3 ;
			RECT 220.477 38.363 220.677 38.461 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 42.395 220.677 42.493 ;
			LAYER M2 ;
			RECT 220.477 42.395 220.677 42.493 ;
			LAYER M3 ;
			RECT 220.477 42.395 220.677 42.493 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 46.427 220.677 46.525 ;
			LAYER M2 ;
			RECT 220.477 46.427 220.677 46.525 ;
			LAYER M3 ;
			RECT 220.477 46.427 220.677 46.525 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 50.459 220.677 50.557 ;
			LAYER M2 ;
			RECT 220.477 50.459 220.677 50.557 ;
			LAYER M3 ;
			RECT 220.477 50.459 220.677 50.557 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 54.491 220.677 54.589 ;
			LAYER M2 ;
			RECT 220.477 54.491 220.677 54.589 ;
			LAYER M3 ;
			RECT 220.477 54.491 220.677 54.589 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 57.515 220.677 57.613 ;
			LAYER M2 ;
			RECT 220.477 57.515 220.677 57.613 ;
			LAYER M3 ;
			RECT 220.477 57.515 220.677 57.613 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 59.531 220.677 59.629 ;
			LAYER M2 ;
			RECT 220.477 59.531 220.677 59.629 ;
			LAYER M3 ;
			RECT 220.477 59.531 220.677 59.629 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 83.299 220.677 83.397 ;
			LAYER M2 ;
			RECT 220.477 83.299 220.677 83.397 ;
			LAYER M3 ;
			RECT 220.477 83.299 220.677 83.397 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 85.355 220.677 85.453 ;
			LAYER M2 ;
			RECT 220.477 85.355 220.677 85.453 ;
			LAYER M3 ;
			RECT 220.477 85.355 220.677 85.453 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 88.379 220.677 88.477 ;
			LAYER M2 ;
			RECT 220.477 88.379 220.677 88.477 ;
			LAYER M3 ;
			RECT 220.477 88.379 220.677 88.477 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 92.411 220.677 92.509 ;
			LAYER M2 ;
			RECT 220.477 92.411 220.677 92.509 ;
			LAYER M3 ;
			RECT 220.477 92.411 220.677 92.509 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 96.443 220.677 96.541 ;
			LAYER M2 ;
			RECT 220.477 96.443 220.677 96.541 ;
			LAYER M3 ;
			RECT 220.477 96.443 220.677 96.541 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 100.475 220.677 100.573 ;
			LAYER M2 ;
			RECT 220.477 100.475 220.677 100.573 ;
			LAYER M3 ;
			RECT 220.477 100.475 220.677 100.573 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 104.507 220.677 104.605 ;
			LAYER M2 ;
			RECT 220.477 104.507 220.677 104.605 ;
			LAYER M3 ;
			RECT 220.477 104.507 220.677 104.605 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 108.539 220.677 108.637 ;
			LAYER M2 ;
			RECT 220.477 108.539 220.677 108.637 ;
			LAYER M3 ;
			RECT 220.477 108.539 220.677 108.637 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 112.571 220.677 112.669 ;
			LAYER M2 ;
			RECT 220.477 112.571 220.677 112.669 ;
			LAYER M3 ;
			RECT 220.477 112.571 220.677 112.669 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 116.603 220.677 116.701 ;
			LAYER M2 ;
			RECT 220.477 116.603 220.677 116.701 ;
			LAYER M3 ;
			RECT 220.477 116.603 220.677 116.701 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 120.635 220.677 120.733 ;
			LAYER M2 ;
			RECT 220.477 120.635 220.677 120.733 ;
			LAYER M3 ;
			RECT 220.477 120.635 220.677 120.733 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 124.667 220.677 124.765 ;
			LAYER M2 ;
			RECT 220.477 124.667 220.677 124.765 ;
			LAYER M3 ;
			RECT 220.477 124.667 220.677 124.765 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 128.699 220.677 128.797 ;
			LAYER M2 ;
			RECT 220.477 128.699 220.677 128.797 ;
			LAYER M3 ;
			RECT 220.477 128.699 220.677 128.797 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 132.731 220.677 132.829 ;
			LAYER M2 ;
			RECT 220.477 132.731 220.677 132.829 ;
			LAYER M3 ;
			RECT 220.477 132.731 220.677 132.829 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 136.763 220.677 136.861 ;
			LAYER M2 ;
			RECT 220.477 136.763 220.677 136.861 ;
			LAYER M3 ;
			RECT 220.477 136.763 220.677 136.861 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 140.795 220.677 140.893 ;
			LAYER M2 ;
			RECT 220.477 140.795 220.677 140.893 ;
			LAYER M3 ;
			RECT 220.477 140.795 220.677 140.893 ;
		END
		ANTENNADIFFAREA 0.048400 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.153840 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.007320 LAYER VIA1 ;
		ANTENNADIFFAREA 0.048400 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.332160 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNADIFFAREA 0.048400 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.682440 LAYER M3 ;
	END Q[31]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 67.367 220.677 67.465 ;
			LAYER M2 ;
			RECT 220.477 67.367 220.677 67.465 ;
			LAYER M3 ;
			RECT 220.477 67.367 220.677 67.465 ;
		END
		ANTENNAGATEAREA 0.009400 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.440160 LAYER M1 ;
		ANTENNAMAXAREACAR 19.138000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009400 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.566120 LAYER M2 ;
		ANTENNAMAXAREACAR 731.670000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009400 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.406520 LAYER M3 ;
		ANTENNAMAXAREACAR 792.931000 LAYER M3 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 68.787 220.677 68.885 ;
			LAYER M2 ;
			RECT 220.477 68.787 220.677 68.885 ;
			LAYER M3 ;
			RECT 220.477 68.787 220.677 68.885 ;
		END
		ANTENNAGATEAREA 0.009400 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.440160 LAYER M1 ;
		ANTENNAMAXAREACAR 19.138000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.012240 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.059360 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009400 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.566120 LAYER M2 ;
		ANTENNAMAXAREACAR 731.670000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.011040 LAYER VIA2 ;
		ANTENNAMAXAREACAR 2.383440 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009400 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.406520 LAYER M3 ;
		ANTENNAMAXAREACAR 792.931000 LAYER M3 ;
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 2.028 220.557 2.148 ;
			LAYER M4 ;
			RECT 0.120 2.776 220.557 2.896 ;
			LAYER M4 ;
			RECT 0.120 3.056 220.557 3.176 ;
			LAYER M4 ;
			RECT 0.120 3.804 220.557 3.924 ;
			LAYER M4 ;
			RECT 0.120 4.224 220.557 4.344 ;
			LAYER M4 ;
			RECT 0.120 6.060 220.557 6.180 ;
			LAYER M4 ;
			RECT 0.120 6.808 220.557 6.928 ;
			LAYER M4 ;
			RECT 0.120 7.088 220.557 7.208 ;
			LAYER M4 ;
			RECT 0.120 7.836 220.557 7.956 ;
			LAYER M4 ;
			RECT 0.120 8.256 220.557 8.376 ;
			LAYER M4 ;
			RECT 0.120 10.092 220.557 10.212 ;
			LAYER M4 ;
			RECT 0.120 10.840 220.557 10.960 ;
			LAYER M4 ;
			RECT 0.120 11.120 220.557 11.240 ;
			LAYER M4 ;
			RECT 0.120 11.868 220.557 11.988 ;
			LAYER M4 ;
			RECT 0.120 12.288 220.557 12.408 ;
			LAYER M4 ;
			RECT 0.120 14.124 220.557 14.244 ;
			LAYER M4 ;
			RECT 0.120 14.872 220.557 14.992 ;
			LAYER M4 ;
			RECT 0.120 15.152 220.557 15.272 ;
			LAYER M4 ;
			RECT 0.120 15.900 220.557 16.020 ;
			LAYER M4 ;
			RECT 0.120 16.320 220.557 16.440 ;
			LAYER M4 ;
			RECT 0.120 18.156 220.557 18.276 ;
			LAYER M4 ;
			RECT 0.120 18.904 220.557 19.024 ;
			LAYER M4 ;
			RECT 0.120 19.184 220.557 19.304 ;
			LAYER M4 ;
			RECT 0.120 19.932 220.557 20.052 ;
			LAYER M4 ;
			RECT 0.120 20.352 220.557 20.472 ;
			LAYER M4 ;
			RECT 0.120 22.188 220.557 22.308 ;
			LAYER M4 ;
			RECT 0.120 22.936 220.557 23.056 ;
			LAYER M4 ;
			RECT 0.120 23.216 220.557 23.336 ;
			LAYER M4 ;
			RECT 0.120 23.964 220.557 24.084 ;
			LAYER M4 ;
			RECT 0.120 24.384 220.557 24.504 ;
			LAYER M4 ;
			RECT 0.120 26.220 220.557 26.340 ;
			LAYER M4 ;
			RECT 0.120 26.968 220.557 27.088 ;
			LAYER M4 ;
			RECT 0.120 27.248 220.557 27.368 ;
			LAYER M4 ;
			RECT 0.120 27.996 220.557 28.116 ;
			LAYER M4 ;
			RECT 0.120 28.416 220.557 28.536 ;
			LAYER M4 ;
			RECT 0.120 30.252 220.557 30.372 ;
			LAYER M4 ;
			RECT 0.120 31.000 220.557 31.120 ;
			LAYER M4 ;
			RECT 0.120 31.280 220.557 31.400 ;
			LAYER M4 ;
			RECT 0.120 32.028 220.557 32.148 ;
			LAYER M4 ;
			RECT 0.120 32.448 220.557 32.568 ;
			LAYER M4 ;
			RECT 0.120 34.284 220.557 34.404 ;
			LAYER M4 ;
			RECT 0.120 35.032 220.557 35.152 ;
			LAYER M4 ;
			RECT 0.120 35.312 220.557 35.432 ;
			LAYER M4 ;
			RECT 0.120 36.060 220.557 36.180 ;
			LAYER M4 ;
			RECT 0.120 36.480 220.557 36.600 ;
			LAYER M4 ;
			RECT 0.120 38.316 220.557 38.436 ;
			LAYER M4 ;
			RECT 0.120 39.064 220.557 39.184 ;
			LAYER M4 ;
			RECT 0.120 39.344 220.557 39.464 ;
			LAYER M4 ;
			RECT 0.120 40.092 220.557 40.212 ;
			LAYER M4 ;
			RECT 0.120 40.512 220.557 40.632 ;
			LAYER M4 ;
			RECT 0.120 42.348 220.557 42.468 ;
			LAYER M4 ;
			RECT 0.120 43.096 220.557 43.216 ;
			LAYER M4 ;
			RECT 0.120 43.376 220.557 43.496 ;
			LAYER M4 ;
			RECT 0.120 44.124 220.557 44.244 ;
			LAYER M4 ;
			RECT 0.120 44.544 220.557 44.664 ;
			LAYER M4 ;
			RECT 0.120 46.380 220.557 46.500 ;
			LAYER M4 ;
			RECT 0.120 47.128 220.557 47.248 ;
			LAYER M4 ;
			RECT 0.120 47.408 220.557 47.528 ;
			LAYER M4 ;
			RECT 0.120 48.156 220.557 48.276 ;
			LAYER M4 ;
			RECT 0.120 48.576 220.557 48.696 ;
			LAYER M4 ;
			RECT 0.120 50.412 220.557 50.532 ;
			LAYER M4 ;
			RECT 0.120 51.160 220.557 51.280 ;
			LAYER M4 ;
			RECT 0.120 51.440 220.557 51.560 ;
			LAYER M4 ;
			RECT 0.120 52.188 220.557 52.308 ;
			LAYER M4 ;
			RECT 0.120 52.608 220.557 52.728 ;
			LAYER M4 ;
			RECT 0.120 54.444 220.557 54.564 ;
			LAYER M4 ;
			RECT 0.120 55.192 220.557 55.312 ;
			LAYER M4 ;
			RECT 0.120 55.472 220.557 55.592 ;
			LAYER M4 ;
			RECT 0.120 56.220 220.557 56.340 ;
			LAYER M4 ;
			RECT 0.120 56.640 220.557 56.760 ;
			LAYER M4 ;
			RECT 0.120 58.476 220.557 58.596 ;
			LAYER M4 ;
			RECT 0.120 59.224 220.557 59.344 ;
			LAYER M4 ;
			RECT 0.120 59.504 220.557 59.624 ;
			LAYER M4 ;
			RECT 0.120 60.252 220.557 60.372 ;
			LAYER M4 ;
			RECT 0.120 60.672 220.557 60.792 ;
			LAYER M4 ;
			RECT 0.120 62.508 220.557 62.628 ;
			LAYER M4 ;
			RECT 0.120 63.256 220.557 63.376 ;
			LAYER M4 ;
			RECT 0.120 63.536 220.557 63.656 ;
			LAYER M4 ;
			RECT 0.120 64.284 220.557 64.404 ;
			LAYER M4 ;
			RECT 0.120 64.704 220.557 64.824 ;
			LAYER M4 ;
			RECT 0.120 66.676 220.557 66.796 ;
			LAYER M4 ;
			RECT 0.120 68.656 220.557 68.776 ;
			LAYER M4 ;
			RECT 0.120 70.348 220.557 70.468 ;
			LAYER M4 ;
			RECT 0.120 72.436 220.557 72.556 ;
			LAYER M4 ;
			RECT 0.120 74.260 220.557 74.380 ;
			LAYER M4 ;
			RECT 0.120 76.036 220.557 76.156 ;
			LAYER M4 ;
			RECT 0.120 77.836 220.557 77.956 ;
			LAYER M4 ;
			RECT 0.120 80.268 220.557 80.388 ;
			LAYER M4 ;
			RECT 0.120 81.016 220.557 81.136 ;
			LAYER M4 ;
			RECT 0.120 81.296 220.557 81.416 ;
			LAYER M4 ;
			RECT 0.120 82.044 220.557 82.164 ;
			LAYER M4 ;
			RECT 0.120 82.464 220.557 82.584 ;
			LAYER M4 ;
			RECT 0.120 84.300 220.557 84.420 ;
			LAYER M4 ;
			RECT 0.120 85.048 220.557 85.168 ;
			LAYER M4 ;
			RECT 0.120 85.328 220.557 85.448 ;
			LAYER M4 ;
			RECT 0.120 86.076 220.557 86.196 ;
			LAYER M4 ;
			RECT 0.120 86.496 220.557 86.616 ;
			LAYER M4 ;
			RECT 0.120 88.332 220.557 88.452 ;
			LAYER M4 ;
			RECT 0.120 89.080 220.557 89.200 ;
			LAYER M4 ;
			RECT 0.120 89.360 220.557 89.480 ;
			LAYER M4 ;
			RECT 0.120 90.108 220.557 90.228 ;
			LAYER M4 ;
			RECT 0.120 90.528 220.557 90.648 ;
			LAYER M4 ;
			RECT 0.120 92.364 220.557 92.484 ;
			LAYER M4 ;
			RECT 0.120 93.112 220.557 93.232 ;
			LAYER M4 ;
			RECT 0.120 93.392 220.557 93.512 ;
			LAYER M4 ;
			RECT 0.120 94.140 220.557 94.260 ;
			LAYER M4 ;
			RECT 0.120 94.560 220.557 94.680 ;
			LAYER M4 ;
			RECT 0.120 96.396 220.557 96.516 ;
			LAYER M4 ;
			RECT 0.120 97.144 220.557 97.264 ;
			LAYER M4 ;
			RECT 0.120 97.424 220.557 97.544 ;
			LAYER M4 ;
			RECT 0.120 98.172 220.557 98.292 ;
			LAYER M4 ;
			RECT 0.120 98.592 220.557 98.712 ;
			LAYER M4 ;
			RECT 0.120 100.428 220.557 100.548 ;
			LAYER M4 ;
			RECT 0.120 101.176 220.557 101.296 ;
			LAYER M4 ;
			RECT 0.120 101.456 220.557 101.576 ;
			LAYER M4 ;
			RECT 0.120 102.204 220.557 102.324 ;
			LAYER M4 ;
			RECT 0.120 102.624 220.557 102.744 ;
			LAYER M4 ;
			RECT 0.120 104.460 220.557 104.580 ;
			LAYER M4 ;
			RECT 0.120 105.208 220.557 105.328 ;
			LAYER M4 ;
			RECT 0.120 105.488 220.557 105.608 ;
			LAYER M4 ;
			RECT 0.120 106.236 220.557 106.356 ;
			LAYER M4 ;
			RECT 0.120 106.656 220.557 106.776 ;
			LAYER M4 ;
			RECT 0.120 108.492 220.557 108.612 ;
			LAYER M4 ;
			RECT 0.120 109.240 220.557 109.360 ;
			LAYER M4 ;
			RECT 0.120 109.520 220.557 109.640 ;
			LAYER M4 ;
			RECT 0.120 110.268 220.557 110.388 ;
			LAYER M4 ;
			RECT 0.120 110.688 220.557 110.808 ;
			LAYER M4 ;
			RECT 0.120 112.524 220.557 112.644 ;
			LAYER M4 ;
			RECT 0.120 113.272 220.557 113.392 ;
			LAYER M4 ;
			RECT 0.120 113.552 220.557 113.672 ;
			LAYER M4 ;
			RECT 0.120 114.300 220.557 114.420 ;
			LAYER M4 ;
			RECT 0.120 114.720 220.557 114.840 ;
			LAYER M4 ;
			RECT 0.120 116.556 220.557 116.676 ;
			LAYER M4 ;
			RECT 0.120 117.304 220.557 117.424 ;
			LAYER M4 ;
			RECT 0.120 117.584 220.557 117.704 ;
			LAYER M4 ;
			RECT 0.120 118.332 220.557 118.452 ;
			LAYER M4 ;
			RECT 0.120 118.752 220.557 118.872 ;
			LAYER M4 ;
			RECT 0.120 120.588 220.557 120.708 ;
			LAYER M4 ;
			RECT 0.120 121.336 220.557 121.456 ;
			LAYER M4 ;
			RECT 0.120 121.616 220.557 121.736 ;
			LAYER M4 ;
			RECT 0.120 122.364 220.557 122.484 ;
			LAYER M4 ;
			RECT 0.120 122.784 220.557 122.904 ;
			LAYER M4 ;
			RECT 0.120 124.620 220.557 124.740 ;
			LAYER M4 ;
			RECT 0.120 125.368 220.557 125.488 ;
			LAYER M4 ;
			RECT 0.120 125.648 220.557 125.768 ;
			LAYER M4 ;
			RECT 0.120 126.396 220.557 126.516 ;
			LAYER M4 ;
			RECT 0.120 126.816 220.557 126.936 ;
			LAYER M4 ;
			RECT 0.120 128.652 220.557 128.772 ;
			LAYER M4 ;
			RECT 0.120 129.400 220.557 129.520 ;
			LAYER M4 ;
			RECT 0.120 129.680 220.557 129.800 ;
			LAYER M4 ;
			RECT 0.120 130.428 220.557 130.548 ;
			LAYER M4 ;
			RECT 0.120 130.848 220.557 130.968 ;
			LAYER M4 ;
			RECT 0.120 132.684 220.557 132.804 ;
			LAYER M4 ;
			RECT 0.120 133.432 220.557 133.552 ;
			LAYER M4 ;
			RECT 0.120 133.712 220.557 133.832 ;
			LAYER M4 ;
			RECT 0.120 134.460 220.557 134.580 ;
			LAYER M4 ;
			RECT 0.120 134.880 220.557 135.000 ;
			LAYER M4 ;
			RECT 0.120 136.716 220.557 136.836 ;
			LAYER M4 ;
			RECT 0.120 137.464 220.557 137.584 ;
			LAYER M4 ;
			RECT 0.120 137.744 220.557 137.864 ;
			LAYER M4 ;
			RECT 0.120 138.492 220.557 138.612 ;
			LAYER M4 ;
			RECT 0.120 138.912 220.557 139.032 ;
			LAYER M4 ;
			RECT 0.120 140.748 220.557 140.868 ;
			LAYER M4 ;
			RECT 0.120 141.496 220.557 141.616 ;
			LAYER M4 ;
			RECT 0.120 141.776 220.557 141.896 ;
			LAYER M4 ;
			RECT 0.120 142.524 220.557 142.644 ;
			LAYER M4 ;
			RECT 0.120 142.944 220.557 143.064 ;
			LAYER M4 ;
			RECT 215.557 68.416 220.557 68.536 ;
			LAYER M4 ;
			RECT 215.557 70.108 220.557 70.228 ;
			LAYER M4 ;
			RECT 215.557 74.500 220.557 74.620 ;
			LAYER M4 ;
			RECT 215.557 76.276 220.557 76.396 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 0.900 220.557 1.020 ;
			LAYER M4 ;
			RECT 0.120 1.608 220.557 1.728 ;
			LAYER M4 ;
			RECT 0.120 2.531 220.557 2.651 ;
			LAYER M4 ;
			RECT 0.120 3.301 220.557 3.421 ;
			LAYER M4 ;
			RECT 0.120 4.932 220.557 5.052 ;
			LAYER M4 ;
			RECT 0.120 5.640 220.557 5.760 ;
			LAYER M4 ;
			RECT 0.120 6.563 220.557 6.683 ;
			LAYER M4 ;
			RECT 0.120 7.333 220.557 7.453 ;
			LAYER M4 ;
			RECT 0.120 8.964 220.557 9.084 ;
			LAYER M4 ;
			RECT 0.120 9.672 220.557 9.792 ;
			LAYER M4 ;
			RECT 0.120 10.595 220.557 10.715 ;
			LAYER M4 ;
			RECT 0.120 11.365 220.557 11.485 ;
			LAYER M4 ;
			RECT 0.120 12.996 220.557 13.116 ;
			LAYER M4 ;
			RECT 0.120 13.704 220.557 13.824 ;
			LAYER M4 ;
			RECT 0.120 14.627 220.557 14.747 ;
			LAYER M4 ;
			RECT 0.120 15.397 220.557 15.517 ;
			LAYER M4 ;
			RECT 0.120 17.028 220.557 17.148 ;
			LAYER M4 ;
			RECT 0.120 17.736 220.557 17.856 ;
			LAYER M4 ;
			RECT 0.120 18.659 220.557 18.779 ;
			LAYER M4 ;
			RECT 0.120 19.429 220.557 19.549 ;
			LAYER M4 ;
			RECT 0.120 21.060 220.557 21.180 ;
			LAYER M4 ;
			RECT 0.120 21.768 220.557 21.888 ;
			LAYER M4 ;
			RECT 0.120 22.691 220.557 22.811 ;
			LAYER M4 ;
			RECT 0.120 23.461 220.557 23.581 ;
			LAYER M4 ;
			RECT 0.120 25.092 220.557 25.212 ;
			LAYER M4 ;
			RECT 0.120 25.800 220.557 25.920 ;
			LAYER M4 ;
			RECT 0.120 26.723 220.557 26.843 ;
			LAYER M4 ;
			RECT 0.120 27.493 220.557 27.613 ;
			LAYER M4 ;
			RECT 0.120 29.124 220.557 29.244 ;
			LAYER M4 ;
			RECT 0.120 29.832 220.557 29.952 ;
			LAYER M4 ;
			RECT 0.120 30.755 220.557 30.875 ;
			LAYER M4 ;
			RECT 0.120 31.525 220.557 31.645 ;
			LAYER M4 ;
			RECT 0.120 33.156 220.557 33.276 ;
			LAYER M4 ;
			RECT 0.120 33.864 220.557 33.984 ;
			LAYER M4 ;
			RECT 0.120 34.787 220.557 34.907 ;
			LAYER M4 ;
			RECT 0.120 35.557 220.557 35.677 ;
			LAYER M4 ;
			RECT 0.120 37.188 220.557 37.308 ;
			LAYER M4 ;
			RECT 0.120 37.896 220.557 38.016 ;
			LAYER M4 ;
			RECT 0.120 38.819 220.557 38.939 ;
			LAYER M4 ;
			RECT 0.120 39.589 220.557 39.709 ;
			LAYER M4 ;
			RECT 0.120 41.220 220.557 41.340 ;
			LAYER M4 ;
			RECT 0.120 41.928 220.557 42.048 ;
			LAYER M4 ;
			RECT 0.120 42.851 220.557 42.971 ;
			LAYER M4 ;
			RECT 0.120 43.621 220.557 43.741 ;
			LAYER M4 ;
			RECT 0.120 45.252 220.557 45.372 ;
			LAYER M4 ;
			RECT 0.120 45.960 220.557 46.080 ;
			LAYER M4 ;
			RECT 0.120 46.883 220.557 47.003 ;
			LAYER M4 ;
			RECT 0.120 47.653 220.557 47.773 ;
			LAYER M4 ;
			RECT 0.120 49.284 220.557 49.404 ;
			LAYER M4 ;
			RECT 0.120 49.992 220.557 50.112 ;
			LAYER M4 ;
			RECT 0.120 50.915 220.557 51.035 ;
			LAYER M4 ;
			RECT 0.120 51.685 220.557 51.805 ;
			LAYER M4 ;
			RECT 0.120 53.316 220.557 53.436 ;
			LAYER M4 ;
			RECT 0.120 54.024 220.557 54.144 ;
			LAYER M4 ;
			RECT 0.120 54.947 220.557 55.067 ;
			LAYER M4 ;
			RECT 0.120 55.717 220.557 55.837 ;
			LAYER M4 ;
			RECT 0.120 57.348 220.557 57.468 ;
			LAYER M4 ;
			RECT 0.120 58.056 220.557 58.176 ;
			LAYER M4 ;
			RECT 0.120 58.979 220.557 59.099 ;
			LAYER M4 ;
			RECT 0.120 59.749 220.557 59.869 ;
			LAYER M4 ;
			RECT 0.120 61.380 220.557 61.500 ;
			LAYER M4 ;
			RECT 0.120 62.088 220.557 62.208 ;
			LAYER M4 ;
			RECT 0.120 63.011 220.557 63.131 ;
			LAYER M4 ;
			RECT 0.120 63.781 220.557 63.901 ;
			LAYER M4 ;
			RECT 0.120 65.412 220.557 65.532 ;
			LAYER M4 ;
			RECT 0.120 68.896 220.557 69.016 ;
			LAYER M4 ;
			RECT 0.120 70.588 220.557 70.708 ;
			LAYER M4 ;
			RECT 0.120 74.020 220.557 74.140 ;
			LAYER M4 ;
			RECT 0.120 75.796 220.557 75.916 ;
			LAYER M4 ;
			RECT 0.120 79.140 220.557 79.260 ;
			LAYER M4 ;
			RECT 0.120 79.848 220.557 79.968 ;
			LAYER M4 ;
			RECT 0.120 80.771 220.557 80.891 ;
			LAYER M4 ;
			RECT 0.120 81.541 220.557 81.661 ;
			LAYER M4 ;
			RECT 0.120 83.172 220.557 83.292 ;
			LAYER M4 ;
			RECT 0.120 83.880 220.557 84.000 ;
			LAYER M4 ;
			RECT 0.120 84.803 220.557 84.923 ;
			LAYER M4 ;
			RECT 0.120 85.573 220.557 85.693 ;
			LAYER M4 ;
			RECT 0.120 87.204 220.557 87.324 ;
			LAYER M4 ;
			RECT 0.120 87.912 220.557 88.032 ;
			LAYER M4 ;
			RECT 0.120 88.835 220.557 88.955 ;
			LAYER M4 ;
			RECT 0.120 89.605 220.557 89.725 ;
			LAYER M4 ;
			RECT 0.120 91.236 220.557 91.356 ;
			LAYER M4 ;
			RECT 0.120 91.944 220.557 92.064 ;
			LAYER M4 ;
			RECT 0.120 92.867 220.557 92.987 ;
			LAYER M4 ;
			RECT 0.120 93.637 220.557 93.757 ;
			LAYER M4 ;
			RECT 0.120 95.268 220.557 95.388 ;
			LAYER M4 ;
			RECT 0.120 95.976 220.557 96.096 ;
			LAYER M4 ;
			RECT 0.120 96.899 220.557 97.019 ;
			LAYER M4 ;
			RECT 0.120 97.669 220.557 97.789 ;
			LAYER M4 ;
			RECT 0.120 99.300 220.557 99.420 ;
			LAYER M4 ;
			RECT 0.120 100.008 220.557 100.128 ;
			LAYER M4 ;
			RECT 0.120 100.931 220.557 101.051 ;
			LAYER M4 ;
			RECT 0.120 101.701 220.557 101.821 ;
			LAYER M4 ;
			RECT 0.120 103.332 220.557 103.452 ;
			LAYER M4 ;
			RECT 0.120 104.040 220.557 104.160 ;
			LAYER M4 ;
			RECT 0.120 104.963 220.557 105.083 ;
			LAYER M4 ;
			RECT 0.120 105.733 220.557 105.853 ;
			LAYER M4 ;
			RECT 0.120 107.364 220.557 107.484 ;
			LAYER M4 ;
			RECT 0.120 108.072 220.557 108.192 ;
			LAYER M4 ;
			RECT 0.120 108.995 220.557 109.115 ;
			LAYER M4 ;
			RECT 0.120 109.765 220.557 109.885 ;
			LAYER M4 ;
			RECT 0.120 111.396 220.557 111.516 ;
			LAYER M4 ;
			RECT 0.120 112.104 220.557 112.224 ;
			LAYER M4 ;
			RECT 0.120 113.027 220.557 113.147 ;
			LAYER M4 ;
			RECT 0.120 113.797 220.557 113.917 ;
			LAYER M4 ;
			RECT 0.120 115.428 220.557 115.548 ;
			LAYER M4 ;
			RECT 0.120 116.136 220.557 116.256 ;
			LAYER M4 ;
			RECT 0.120 117.059 220.557 117.179 ;
			LAYER M4 ;
			RECT 0.120 117.829 220.557 117.949 ;
			LAYER M4 ;
			RECT 0.120 119.460 220.557 119.580 ;
			LAYER M4 ;
			RECT 0.120 120.168 220.557 120.288 ;
			LAYER M4 ;
			RECT 0.120 121.091 220.557 121.211 ;
			LAYER M4 ;
			RECT 0.120 121.861 220.557 121.981 ;
			LAYER M4 ;
			RECT 0.120 123.492 220.557 123.612 ;
			LAYER M4 ;
			RECT 0.120 124.200 220.557 124.320 ;
			LAYER M4 ;
			RECT 0.120 125.123 220.557 125.243 ;
			LAYER M4 ;
			RECT 0.120 125.893 220.557 126.013 ;
			LAYER M4 ;
			RECT 0.120 127.524 220.557 127.644 ;
			LAYER M4 ;
			RECT 0.120 128.232 220.557 128.352 ;
			LAYER M4 ;
			RECT 0.120 129.155 220.557 129.275 ;
			LAYER M4 ;
			RECT 0.120 129.925 220.557 130.045 ;
			LAYER M4 ;
			RECT 0.120 131.556 220.557 131.676 ;
			LAYER M4 ;
			RECT 0.120 132.264 220.557 132.384 ;
			LAYER M4 ;
			RECT 0.120 133.187 220.557 133.307 ;
			LAYER M4 ;
			RECT 0.120 133.957 220.557 134.077 ;
			LAYER M4 ;
			RECT 0.120 135.588 220.557 135.708 ;
			LAYER M4 ;
			RECT 0.120 136.296 220.557 136.416 ;
			LAYER M4 ;
			RECT 0.120 137.219 220.557 137.339 ;
			LAYER M4 ;
			RECT 0.120 137.989 220.557 138.109 ;
			LAYER M4 ;
			RECT 0.120 139.620 220.557 139.740 ;
			LAYER M4 ;
			RECT 0.120 140.328 220.557 140.448 ;
			LAYER M4 ;
			RECT 0.120 141.251 220.557 141.371 ;
			LAYER M4 ;
			RECT 0.120 142.021 220.557 142.141 ;
			LAYER M4 ;
			RECT 0.120 143.652 220.557 143.772 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 68.549 220.677 68.647 ;
			LAYER M2 ;
			RECT 220.477 68.549 220.677 68.647 ;
			LAYER M3 ;
			RECT 220.477 68.549 220.677 68.647 ;
		END
		ANTENNAGATEAREA 0.006200 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.142800 LAYER M1 ;
		ANTENNAMAXAREACAR 12.155900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.004920 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.199440 LAYER VIA1 ;
		ANTENNAGATEAREA 0.006200 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.088800 LAYER M2 ;
		ANTENNAMAXAREACAR 14.912300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006120 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.399000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.006200 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085680 LAYER M3 ;
		ANTENNAMAXAREACAR 27.095000 LAYER M3 ;
	END WEB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 69.025 220.677 69.123 ;
			LAYER M2 ;
			RECT 220.477 69.025 220.677 69.123 ;
			LAYER M3 ;
			RECT 220.477 69.025 220.677 69.123 ;
		END
		ANTENNAGATEAREA 0.007100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.280320 LAYER M1 ;
		ANTENNAMAXAREACAR 12.244400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.172560 LAYER VIA1 ;
		ANTENNAGATEAREA 0.007100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.145040 LAYER M2 ;
		ANTENNAMAXAREACAR 77.595500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.018480 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.345120 LAYER VIA2 ;
		ANTENNAGATEAREA 0.007100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.209360 LAYER M3 ;
		ANTENNAMAXAREACAR 211.858000 LAYER M3 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 220.477 70.745 220.677 70.843 ;
			LAYER M2 ;
			RECT 220.477 70.745 220.677 70.843 ;
			LAYER M3 ;
			RECT 220.477 70.745 220.677 70.843 ;
		END
		ANTENNAGATEAREA 0.007100 LAYER M1 ;
		ANTENNADIFFAREA 0.008100 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.280320 LAYER M1 ;
		ANTENNAMAXAREACAR 12.244400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.008640 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.172560 LAYER VIA1 ;
		ANTENNAGATEAREA 0.007100 LAYER M2 ;
		ANTENNADIFFAREA 0.008100 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.145040 LAYER M2 ;
		ANTENNAMAXAREACAR 77.595500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.018480 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.345120 LAYER VIA2 ;
		ANTENNAGATEAREA 0.007100 LAYER M3 ;
		ANTENNADIFFAREA 0.008100 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.209360 LAYER M3 ;
		ANTENNAMAXAREACAR 211.858000 LAYER M3 ;
	END WTSEL[1]

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 220.677 144.672 ;
		LAYER M2 ;
		RECT 0.000 0.000 220.677 144.672 ;
		LAYER M3 ;
		RECT 0.000 0.000 220.677 144.672 ;
		LAYER M4 ;
		RECT 0.702 69.087 209.653 69.185 ;
		LAYER M4 ;
		RECT 0.702 69.547 213.881 69.645 ;
		LAYER M4 ;
		RECT 0.750 2.179 212.089 2.277 ;
		LAYER M4 ;
		RECT 0.750 3.675 212.089 3.773 ;
		LAYER M4 ;
		RECT 0.750 6.211 212.089 6.309 ;
		LAYER M4 ;
		RECT 0.750 7.707 212.089 7.805 ;
		LAYER M4 ;
		RECT 0.750 10.243 212.089 10.341 ;
		LAYER M4 ;
		RECT 0.750 11.739 212.089 11.837 ;
		LAYER M4 ;
		RECT 0.750 14.275 212.089 14.373 ;
		LAYER M4 ;
		RECT 0.750 15.771 212.089 15.869 ;
		LAYER M4 ;
		RECT 0.750 18.307 212.089 18.405 ;
		LAYER M4 ;
		RECT 0.750 19.803 212.089 19.901 ;
		LAYER M4 ;
		RECT 0.750 22.339 212.089 22.437 ;
		LAYER M4 ;
		RECT 0.750 23.835 212.089 23.933 ;
		LAYER M4 ;
		RECT 0.750 26.371 212.089 26.469 ;
		LAYER M4 ;
		RECT 0.750 27.867 212.089 27.965 ;
		LAYER M4 ;
		RECT 0.750 30.403 212.089 30.501 ;
		LAYER M4 ;
		RECT 0.750 31.899 212.089 31.997 ;
		LAYER M4 ;
		RECT 0.750 34.435 212.089 34.533 ;
		LAYER M4 ;
		RECT 0.750 35.931 212.089 36.029 ;
		LAYER M4 ;
		RECT 0.750 38.467 212.089 38.565 ;
		LAYER M4 ;
		RECT 0.750 39.963 212.089 40.061 ;
		LAYER M4 ;
		RECT 0.750 42.499 212.089 42.597 ;
		LAYER M4 ;
		RECT 0.750 43.995 212.089 44.093 ;
		LAYER M4 ;
		RECT 0.750 46.531 212.089 46.629 ;
		LAYER M4 ;
		RECT 0.750 48.027 212.089 48.125 ;
		LAYER M4 ;
		RECT 0.750 50.563 212.089 50.661 ;
		LAYER M4 ;
		RECT 0.750 52.059 212.089 52.157 ;
		LAYER M4 ;
		RECT 0.750 54.595 212.089 54.693 ;
		LAYER M4 ;
		RECT 0.750 56.091 212.089 56.189 ;
		LAYER M4 ;
		RECT 0.750 58.627 208.623 58.725 ;
		LAYER M4 ;
		RECT 0.750 60.123 209.112 60.221 ;
		LAYER M4 ;
		RECT 0.750 62.659 209.859 62.757 ;
		LAYER M4 ;
		RECT 0.750 64.155 209.433 64.253 ;
		LAYER M4 ;
		RECT 0.750 65.673 209.047 65.771 ;
		LAYER M4 ;
		RECT 0.750 65.831 209.157 65.929 ;
		LAYER M4 ;
		RECT 0.750 65.989 209.839 66.087 ;
		LAYER M4 ;
		RECT 0.750 66.147 212.107 66.245 ;
		LAYER M4 ;
		RECT 0.750 66.507 209.425 66.605 ;
		LAYER M4 ;
		RECT 0.750 67.047 212.395 67.145 ;
		LAYER M4 ;
		RECT 0.750 67.227 209.047 67.325 ;
		LAYER M4 ;
		RECT 0.750 67.407 212.485 67.505 ;
		LAYER M4 ;
		RECT 0.750 67.587 209.047 67.685 ;
		LAYER M4 ;
		RECT 0.750 67.767 212.395 67.865 ;
		LAYER M4 ;
		RECT 0.750 67.947 209.157 68.045 ;
		LAYER M4 ;
		RECT 0.750 68.127 212.127 68.225 ;
		LAYER M4 ;
		RECT 0.750 68.307 209.047 68.405 ;
		LAYER M4 ;
		RECT 0.750 70.827 213.297 70.925 ;
		LAYER M4 ;
		RECT 0.750 71.007 212.127 71.105 ;
		LAYER M4 ;
		RECT 0.750 71.187 209.425 71.285 ;
		LAYER M4 ;
		RECT 0.750 71.367 214.421 71.465 ;
		LAYER M4 ;
		RECT 0.750 71.547 215.590 71.645 ;
		LAYER M4 ;
		RECT 0.750 71.727 211.086 71.825 ;
		LAYER M4 ;
		RECT 0.750 71.907 215.501 72.005 ;
		LAYER M4 ;
		RECT 0.750 72.087 211.321 72.185 ;
		LAYER M4 ;
		RECT 0.750 72.745 214.061 72.843 ;
		LAYER M4 ;
		RECT 0.750 72.903 209.047 73.001 ;
		LAYER M4 ;
		RECT 0.750 73.061 213.881 73.159 ;
		LAYER M4 ;
		RECT 0.750 73.219 209.160 73.317 ;
		LAYER M4 ;
		RECT 0.750 73.377 211.321 73.475 ;
		LAYER M4 ;
		RECT 0.750 73.535 211.321 73.633 ;
		LAYER M4 ;
		RECT 0.750 73.693 213.881 73.791 ;
		LAYER M4 ;
		RECT 0.750 73.851 211.321 73.949 ;
		LAYER M4 ;
		RECT 0.750 75.017 214.781 75.115 ;
		LAYER M4 ;
		RECT 0.750 75.175 209.157 75.273 ;
		LAYER M4 ;
		RECT 0.750 75.333 213.881 75.431 ;
		LAYER M4 ;
		RECT 0.750 75.491 211.091 75.589 ;
		LAYER M4 ;
		RECT 0.750 75.649 209.047 75.747 ;
		LAYER M4 ;
		RECT 0.750 76.407 212.127 76.505 ;
		LAYER M4 ;
		RECT 0.750 76.587 209.157 76.685 ;
		LAYER M4 ;
		RECT 0.750 76.767 212.127 76.865 ;
		LAYER M4 ;
		RECT 0.750 76.947 209.047 77.045 ;
		LAYER M4 ;
		RECT 0.750 77.127 212.377 77.225 ;
		LAYER M4 ;
		RECT 0.750 77.307 209.157 77.405 ;
		LAYER M4 ;
		RECT 0.750 77.487 212.127 77.585 ;
		LAYER M4 ;
		RECT 0.750 77.667 209.047 77.765 ;
		LAYER M4 ;
		RECT 0.750 78.567 212.269 78.665 ;
		LAYER M4 ;
		RECT 0.750 80.419 209.087 80.517 ;
		LAYER M4 ;
		RECT 0.750 81.915 209.447 82.013 ;
		LAYER M4 ;
		RECT 0.750 84.451 209.881 84.549 ;
		LAYER M4 ;
		RECT 0.750 85.947 209.097 86.045 ;
		LAYER M4 ;
		RECT 0.750 88.483 212.089 88.581 ;
		LAYER M4 ;
		RECT 0.750 89.979 212.089 90.077 ;
		LAYER M4 ;
		RECT 0.750 92.515 212.089 92.613 ;
		LAYER M4 ;
		RECT 0.750 94.011 212.089 94.109 ;
		LAYER M4 ;
		RECT 0.750 96.547 212.089 96.645 ;
		LAYER M4 ;
		RECT 0.750 98.043 212.089 98.141 ;
		LAYER M4 ;
		RECT 0.750 100.579 212.089 100.677 ;
		LAYER M4 ;
		RECT 0.750 102.075 212.089 102.173 ;
		LAYER M4 ;
		RECT 0.750 104.611 212.089 104.709 ;
		LAYER M4 ;
		RECT 0.750 106.107 212.089 106.205 ;
		LAYER M4 ;
		RECT 0.750 108.643 212.089 108.741 ;
		LAYER M4 ;
		RECT 0.750 110.139 212.089 110.237 ;
		LAYER M4 ;
		RECT 0.750 112.675 212.089 112.773 ;
		LAYER M4 ;
		RECT 0.750 114.171 212.089 114.269 ;
		LAYER M4 ;
		RECT 0.750 116.707 212.089 116.805 ;
		LAYER M4 ;
		RECT 0.750 118.203 212.089 118.301 ;
		LAYER M4 ;
		RECT 0.750 120.739 212.089 120.837 ;
		LAYER M4 ;
		RECT 0.750 122.235 212.089 122.333 ;
		LAYER M4 ;
		RECT 0.750 124.771 212.089 124.869 ;
		LAYER M4 ;
		RECT 0.750 126.267 212.089 126.365 ;
		LAYER M4 ;
		RECT 0.750 128.803 212.089 128.901 ;
		LAYER M4 ;
		RECT 0.750 130.299 212.089 130.397 ;
		LAYER M4 ;
		RECT 0.750 132.835 212.089 132.933 ;
		LAYER M4 ;
		RECT 0.750 134.331 212.089 134.429 ;
		LAYER M4 ;
		RECT 0.750 136.867 212.089 136.965 ;
		LAYER M4 ;
		RECT 0.750 138.363 212.089 138.461 ;
		LAYER M4 ;
		RECT 0.750 140.899 212.089 140.997 ;
		LAYER M4 ;
		RECT 0.750 142.395 212.089 142.493 ;
		LAYER M4 ;
		RECT 48.847 3.207 52.805 3.259 ;
		LAYER M4 ;
		RECT 48.847 3.441 52.805 3.493 ;
		LAYER M4 ;
		RECT 48.847 7.239 52.805 7.291 ;
		LAYER M4 ;
		RECT 48.847 7.473 52.805 7.525 ;
		LAYER M4 ;
		RECT 48.847 11.271 52.805 11.323 ;
		LAYER M4 ;
		RECT 48.847 11.505 52.805 11.557 ;
		LAYER M4 ;
		RECT 48.847 15.303 52.805 15.355 ;
		LAYER M4 ;
		RECT 48.847 15.537 52.805 15.589 ;
		LAYER M4 ;
		RECT 48.847 19.335 52.805 19.387 ;
		LAYER M4 ;
		RECT 48.847 19.569 52.805 19.621 ;
		LAYER M4 ;
		RECT 48.847 23.367 52.805 23.419 ;
		LAYER M4 ;
		RECT 48.847 23.601 52.805 23.653 ;
		LAYER M4 ;
		RECT 48.847 27.399 52.805 27.451 ;
		LAYER M4 ;
		RECT 48.847 27.633 52.805 27.685 ;
		LAYER M4 ;
		RECT 48.847 31.431 52.805 31.483 ;
		LAYER M4 ;
		RECT 48.847 31.665 52.805 31.717 ;
		LAYER M4 ;
		RECT 48.847 35.463 52.805 35.515 ;
		LAYER M4 ;
		RECT 48.847 35.697 52.805 35.749 ;
		LAYER M4 ;
		RECT 48.847 39.495 52.805 39.547 ;
		LAYER M4 ;
		RECT 48.847 39.729 52.805 39.781 ;
		LAYER M4 ;
		RECT 48.847 43.527 52.805 43.579 ;
		LAYER M4 ;
		RECT 48.847 43.761 52.805 43.813 ;
		LAYER M4 ;
		RECT 48.847 47.559 52.805 47.611 ;
		LAYER M4 ;
		RECT 48.847 47.793 52.805 47.845 ;
		LAYER M4 ;
		RECT 48.847 51.591 52.805 51.643 ;
		LAYER M4 ;
		RECT 48.847 51.825 52.805 51.877 ;
		LAYER M4 ;
		RECT 48.847 55.623 52.805 55.675 ;
		LAYER M4 ;
		RECT 48.847 55.857 52.805 55.909 ;
		LAYER M4 ;
		RECT 48.847 59.655 52.805 59.707 ;
		LAYER M4 ;
		RECT 48.847 59.889 52.805 59.941 ;
		LAYER M4 ;
		RECT 48.847 63.687 52.805 63.739 ;
		LAYER M4 ;
		RECT 48.847 63.921 52.805 63.973 ;
		LAYER M4 ;
		RECT 48.847 81.447 52.805 81.499 ;
		LAYER M4 ;
		RECT 48.847 81.681 52.805 81.733 ;
		LAYER M4 ;
		RECT 48.847 85.479 52.805 85.531 ;
		LAYER M4 ;
		RECT 48.847 85.713 52.805 85.765 ;
		LAYER M4 ;
		RECT 48.847 89.511 52.805 89.563 ;
		LAYER M4 ;
		RECT 48.847 89.745 52.805 89.797 ;
		LAYER M4 ;
		RECT 48.847 93.543 52.805 93.595 ;
		LAYER M4 ;
		RECT 48.847 93.777 52.805 93.829 ;
		LAYER M4 ;
		RECT 48.847 97.575 52.805 97.627 ;
		LAYER M4 ;
		RECT 48.847 97.809 52.805 97.861 ;
		LAYER M4 ;
		RECT 48.847 101.607 52.805 101.659 ;
		LAYER M4 ;
		RECT 48.847 101.841 52.805 101.893 ;
		LAYER M4 ;
		RECT 48.847 105.639 52.805 105.691 ;
		LAYER M4 ;
		RECT 48.847 105.873 52.805 105.925 ;
		LAYER M4 ;
		RECT 48.847 109.671 52.805 109.723 ;
		LAYER M4 ;
		RECT 48.847 109.905 52.805 109.957 ;
		LAYER M4 ;
		RECT 48.847 113.703 52.805 113.755 ;
		LAYER M4 ;
		RECT 48.847 113.937 52.805 113.989 ;
		LAYER M4 ;
		RECT 48.847 117.735 52.805 117.787 ;
		LAYER M4 ;
		RECT 48.847 117.969 52.805 118.021 ;
		LAYER M4 ;
		RECT 48.847 121.767 52.805 121.819 ;
		LAYER M4 ;
		RECT 48.847 122.001 52.805 122.053 ;
		LAYER M4 ;
		RECT 48.847 125.799 52.805 125.851 ;
		LAYER M4 ;
		RECT 48.847 126.033 52.805 126.085 ;
		LAYER M4 ;
		RECT 48.847 129.831 52.805 129.883 ;
		LAYER M4 ;
		RECT 48.847 130.065 52.805 130.117 ;
		LAYER M4 ;
		RECT 48.847 133.863 52.805 133.915 ;
		LAYER M4 ;
		RECT 48.847 134.097 52.805 134.149 ;
		LAYER M4 ;
		RECT 48.847 137.895 52.805 137.947 ;
		LAYER M4 ;
		RECT 48.847 138.129 52.805 138.181 ;
		LAYER M4 ;
		RECT 48.847 141.927 52.805 141.979 ;
		LAYER M4 ;
		RECT 48.847 142.161 52.805 142.213 ;
		LAYER M4 ;
		RECT 52.543 2.459 56.501 2.511 ;
		LAYER M4 ;
		RECT 52.543 2.693 56.501 2.745 ;
		LAYER M4 ;
		RECT 52.543 6.491 56.501 6.543 ;
		LAYER M4 ;
		RECT 52.543 6.725 56.501 6.777 ;
		LAYER M4 ;
		RECT 52.543 10.523 56.501 10.575 ;
		LAYER M4 ;
		RECT 52.543 10.757 56.501 10.809 ;
		LAYER M4 ;
		RECT 52.543 14.555 56.501 14.607 ;
		LAYER M4 ;
		RECT 52.543 14.789 56.501 14.841 ;
		LAYER M4 ;
		RECT 52.543 18.587 56.501 18.639 ;
		LAYER M4 ;
		RECT 52.543 18.821 56.501 18.873 ;
		LAYER M4 ;
		RECT 52.543 22.619 56.501 22.671 ;
		LAYER M4 ;
		RECT 52.543 22.853 56.501 22.905 ;
		LAYER M4 ;
		RECT 52.543 26.651 56.501 26.703 ;
		LAYER M4 ;
		RECT 52.543 26.885 56.501 26.937 ;
		LAYER M4 ;
		RECT 52.543 30.683 56.501 30.735 ;
		LAYER M4 ;
		RECT 52.543 30.917 56.501 30.969 ;
		LAYER M4 ;
		RECT 52.543 34.715 56.501 34.767 ;
		LAYER M4 ;
		RECT 52.543 34.949 56.501 35.001 ;
		LAYER M4 ;
		RECT 52.543 38.747 56.501 38.799 ;
		LAYER M4 ;
		RECT 52.543 38.981 56.501 39.033 ;
		LAYER M4 ;
		RECT 52.543 42.779 56.501 42.831 ;
		LAYER M4 ;
		RECT 52.543 43.013 56.501 43.065 ;
		LAYER M4 ;
		RECT 52.543 46.811 56.501 46.863 ;
		LAYER M4 ;
		RECT 52.543 47.045 56.501 47.097 ;
		LAYER M4 ;
		RECT 52.543 50.843 56.501 50.895 ;
		LAYER M4 ;
		RECT 52.543 51.077 56.501 51.129 ;
		LAYER M4 ;
		RECT 52.543 54.875 56.501 54.927 ;
		LAYER M4 ;
		RECT 52.543 55.109 56.501 55.161 ;
		LAYER M4 ;
		RECT 52.543 58.907 56.501 58.959 ;
		LAYER M4 ;
		RECT 52.543 59.141 56.501 59.193 ;
		LAYER M4 ;
		RECT 52.543 62.939 56.501 62.991 ;
		LAYER M4 ;
		RECT 52.543 63.173 56.501 63.225 ;
		LAYER M4 ;
		RECT 52.543 80.699 56.501 80.751 ;
		LAYER M4 ;
		RECT 52.543 80.933 56.501 80.985 ;
		LAYER M4 ;
		RECT 52.543 84.731 56.501 84.783 ;
		LAYER M4 ;
		RECT 52.543 84.965 56.501 85.017 ;
		LAYER M4 ;
		RECT 52.543 88.763 56.501 88.815 ;
		LAYER M4 ;
		RECT 52.543 88.997 56.501 89.049 ;
		LAYER M4 ;
		RECT 52.543 92.795 56.501 92.847 ;
		LAYER M4 ;
		RECT 52.543 93.029 56.501 93.081 ;
		LAYER M4 ;
		RECT 52.543 96.827 56.501 96.879 ;
		LAYER M4 ;
		RECT 52.543 97.061 56.501 97.113 ;
		LAYER M4 ;
		RECT 52.543 100.859 56.501 100.911 ;
		LAYER M4 ;
		RECT 52.543 101.093 56.501 101.145 ;
		LAYER M4 ;
		RECT 52.543 104.891 56.501 104.943 ;
		LAYER M4 ;
		RECT 52.543 105.125 56.501 105.177 ;
		LAYER M4 ;
		RECT 52.543 108.923 56.501 108.975 ;
		LAYER M4 ;
		RECT 52.543 109.157 56.501 109.209 ;
		LAYER M4 ;
		RECT 52.543 112.955 56.501 113.007 ;
		LAYER M4 ;
		RECT 52.543 113.189 56.501 113.241 ;
		LAYER M4 ;
		RECT 52.543 116.987 56.501 117.039 ;
		LAYER M4 ;
		RECT 52.543 117.221 56.501 117.273 ;
		LAYER M4 ;
		RECT 52.543 121.019 56.501 121.071 ;
		LAYER M4 ;
		RECT 52.543 121.253 56.501 121.305 ;
		LAYER M4 ;
		RECT 52.543 125.051 56.501 125.103 ;
		LAYER M4 ;
		RECT 52.543 125.285 56.501 125.337 ;
		LAYER M4 ;
		RECT 52.543 129.083 56.501 129.135 ;
		LAYER M4 ;
		RECT 52.543 129.317 56.501 129.369 ;
		LAYER M4 ;
		RECT 52.543 133.115 56.501 133.167 ;
		LAYER M4 ;
		RECT 52.543 133.349 56.501 133.401 ;
		LAYER M4 ;
		RECT 52.543 137.147 56.501 137.199 ;
		LAYER M4 ;
		RECT 52.543 137.381 56.501 137.433 ;
		LAYER M4 ;
		RECT 52.543 141.179 56.501 141.231 ;
		LAYER M4 ;
		RECT 52.543 141.413 56.501 141.465 ;
		LAYER M4 ;
		RECT 152.287 3.207 156.245 3.259 ;
		LAYER M4 ;
		RECT 152.287 3.441 156.245 3.493 ;
		LAYER M4 ;
		RECT 152.287 7.239 156.245 7.291 ;
		LAYER M4 ;
		RECT 152.287 7.473 156.245 7.525 ;
		LAYER M4 ;
		RECT 152.287 11.271 156.245 11.323 ;
		LAYER M4 ;
		RECT 152.287 11.505 156.245 11.557 ;
		LAYER M4 ;
		RECT 152.287 15.303 156.245 15.355 ;
		LAYER M4 ;
		RECT 152.287 15.537 156.245 15.589 ;
		LAYER M4 ;
		RECT 152.287 19.335 156.245 19.387 ;
		LAYER M4 ;
		RECT 152.287 19.569 156.245 19.621 ;
		LAYER M4 ;
		RECT 152.287 23.367 156.245 23.419 ;
		LAYER M4 ;
		RECT 152.287 23.601 156.245 23.653 ;
		LAYER M4 ;
		RECT 152.287 27.399 156.245 27.451 ;
		LAYER M4 ;
		RECT 152.287 27.633 156.245 27.685 ;
		LAYER M4 ;
		RECT 152.287 31.431 156.245 31.483 ;
		LAYER M4 ;
		RECT 152.287 31.665 156.245 31.717 ;
		LAYER M4 ;
		RECT 152.287 35.463 156.245 35.515 ;
		LAYER M4 ;
		RECT 152.287 35.697 156.245 35.749 ;
		LAYER M4 ;
		RECT 152.287 39.495 156.245 39.547 ;
		LAYER M4 ;
		RECT 152.287 39.729 156.245 39.781 ;
		LAYER M4 ;
		RECT 152.287 43.527 156.245 43.579 ;
		LAYER M4 ;
		RECT 152.287 43.761 156.245 43.813 ;
		LAYER M4 ;
		RECT 152.287 47.559 156.245 47.611 ;
		LAYER M4 ;
		RECT 152.287 47.793 156.245 47.845 ;
		LAYER M4 ;
		RECT 152.287 51.591 156.245 51.643 ;
		LAYER M4 ;
		RECT 152.287 51.825 156.245 51.877 ;
		LAYER M4 ;
		RECT 152.287 55.623 156.245 55.675 ;
		LAYER M4 ;
		RECT 152.287 55.857 156.245 55.909 ;
		LAYER M4 ;
		RECT 152.287 59.655 156.245 59.707 ;
		LAYER M4 ;
		RECT 152.287 59.889 156.245 59.941 ;
		LAYER M4 ;
		RECT 152.287 63.687 156.245 63.739 ;
		LAYER M4 ;
		RECT 152.287 63.921 156.245 63.973 ;
		LAYER M4 ;
		RECT 152.287 81.447 156.245 81.499 ;
		LAYER M4 ;
		RECT 152.287 81.681 156.245 81.733 ;
		LAYER M4 ;
		RECT 152.287 85.479 156.245 85.531 ;
		LAYER M4 ;
		RECT 152.287 85.713 156.245 85.765 ;
		LAYER M4 ;
		RECT 152.287 89.511 156.245 89.563 ;
		LAYER M4 ;
		RECT 152.287 89.745 156.245 89.797 ;
		LAYER M4 ;
		RECT 152.287 93.543 156.245 93.595 ;
		LAYER M4 ;
		RECT 152.287 93.777 156.245 93.829 ;
		LAYER M4 ;
		RECT 152.287 97.575 156.245 97.627 ;
		LAYER M4 ;
		RECT 152.287 97.809 156.245 97.861 ;
		LAYER M4 ;
		RECT 152.287 101.607 156.245 101.659 ;
		LAYER M4 ;
		RECT 152.287 101.841 156.245 101.893 ;
		LAYER M4 ;
		RECT 152.287 105.639 156.245 105.691 ;
		LAYER M4 ;
		RECT 152.287 105.873 156.245 105.925 ;
		LAYER M4 ;
		RECT 152.287 109.671 156.245 109.723 ;
		LAYER M4 ;
		RECT 152.287 109.905 156.245 109.957 ;
		LAYER M4 ;
		RECT 152.287 113.703 156.245 113.755 ;
		LAYER M4 ;
		RECT 152.287 113.937 156.245 113.989 ;
		LAYER M4 ;
		RECT 152.287 117.735 156.245 117.787 ;
		LAYER M4 ;
		RECT 152.287 117.969 156.245 118.021 ;
		LAYER M4 ;
		RECT 152.287 121.767 156.245 121.819 ;
		LAYER M4 ;
		RECT 152.287 122.001 156.245 122.053 ;
		LAYER M4 ;
		RECT 152.287 125.799 156.245 125.851 ;
		LAYER M4 ;
		RECT 152.287 126.033 156.245 126.085 ;
		LAYER M4 ;
		RECT 152.287 129.831 156.245 129.883 ;
		LAYER M4 ;
		RECT 152.287 130.065 156.245 130.117 ;
		LAYER M4 ;
		RECT 152.287 133.863 156.245 133.915 ;
		LAYER M4 ;
		RECT 152.287 134.097 156.245 134.149 ;
		LAYER M4 ;
		RECT 152.287 137.895 156.245 137.947 ;
		LAYER M4 ;
		RECT 152.287 138.129 156.245 138.181 ;
		LAYER M4 ;
		RECT 152.287 141.927 156.245 141.979 ;
		LAYER M4 ;
		RECT 152.287 142.161 156.245 142.213 ;
		LAYER M4 ;
		RECT 155.983 2.459 159.941 2.511 ;
		LAYER M4 ;
		RECT 155.983 2.693 159.941 2.745 ;
		LAYER M4 ;
		RECT 155.983 6.491 159.941 6.543 ;
		LAYER M4 ;
		RECT 155.983 6.725 159.941 6.777 ;
		LAYER M4 ;
		RECT 155.983 10.523 159.941 10.575 ;
		LAYER M4 ;
		RECT 155.983 10.757 159.941 10.809 ;
		LAYER M4 ;
		RECT 155.983 14.555 159.941 14.607 ;
		LAYER M4 ;
		RECT 155.983 14.789 159.941 14.841 ;
		LAYER M4 ;
		RECT 155.983 18.587 159.941 18.639 ;
		LAYER M4 ;
		RECT 155.983 18.821 159.941 18.873 ;
		LAYER M4 ;
		RECT 155.983 22.619 159.941 22.671 ;
		LAYER M4 ;
		RECT 155.983 22.853 159.941 22.905 ;
		LAYER M4 ;
		RECT 155.983 26.651 159.941 26.703 ;
		LAYER M4 ;
		RECT 155.983 26.885 159.941 26.937 ;
		LAYER M4 ;
		RECT 155.983 30.683 159.941 30.735 ;
		LAYER M4 ;
		RECT 155.983 30.917 159.941 30.969 ;
		LAYER M4 ;
		RECT 155.983 34.715 159.941 34.767 ;
		LAYER M4 ;
		RECT 155.983 34.949 159.941 35.001 ;
		LAYER M4 ;
		RECT 155.983 38.747 159.941 38.799 ;
		LAYER M4 ;
		RECT 155.983 38.981 159.941 39.033 ;
		LAYER M4 ;
		RECT 155.983 42.779 159.941 42.831 ;
		LAYER M4 ;
		RECT 155.983 43.013 159.941 43.065 ;
		LAYER M4 ;
		RECT 155.983 46.811 159.941 46.863 ;
		LAYER M4 ;
		RECT 155.983 47.045 159.941 47.097 ;
		LAYER M4 ;
		RECT 155.983 50.843 159.941 50.895 ;
		LAYER M4 ;
		RECT 155.983 51.077 159.941 51.129 ;
		LAYER M4 ;
		RECT 155.983 54.875 159.941 54.927 ;
		LAYER M4 ;
		RECT 155.983 55.109 159.941 55.161 ;
		LAYER M4 ;
		RECT 155.983 58.907 159.941 58.959 ;
		LAYER M4 ;
		RECT 155.983 59.141 159.941 59.193 ;
		LAYER M4 ;
		RECT 155.983 62.939 159.941 62.991 ;
		LAYER M4 ;
		RECT 155.983 63.173 159.941 63.225 ;
		LAYER M4 ;
		RECT 155.983 80.699 159.941 80.751 ;
		LAYER M4 ;
		RECT 155.983 80.933 159.941 80.985 ;
		LAYER M4 ;
		RECT 155.983 84.731 159.941 84.783 ;
		LAYER M4 ;
		RECT 155.983 84.965 159.941 85.017 ;
		LAYER M4 ;
		RECT 155.983 88.763 159.941 88.815 ;
		LAYER M4 ;
		RECT 155.983 88.997 159.941 89.049 ;
		LAYER M4 ;
		RECT 155.983 92.795 159.941 92.847 ;
		LAYER M4 ;
		RECT 155.983 93.029 159.941 93.081 ;
		LAYER M4 ;
		RECT 155.983 96.827 159.941 96.879 ;
		LAYER M4 ;
		RECT 155.983 97.061 159.941 97.113 ;
		LAYER M4 ;
		RECT 155.983 100.859 159.941 100.911 ;
		LAYER M4 ;
		RECT 155.983 101.093 159.941 101.145 ;
		LAYER M4 ;
		RECT 155.983 104.891 159.941 104.943 ;
		LAYER M4 ;
		RECT 155.983 105.125 159.941 105.177 ;
		LAYER M4 ;
		RECT 155.983 108.923 159.941 108.975 ;
		LAYER M4 ;
		RECT 155.983 109.157 159.941 109.209 ;
		LAYER M4 ;
		RECT 155.983 112.955 159.941 113.007 ;
		LAYER M4 ;
		RECT 155.983 113.189 159.941 113.241 ;
		LAYER M4 ;
		RECT 155.983 116.987 159.941 117.039 ;
		LAYER M4 ;
		RECT 155.983 117.221 159.941 117.273 ;
		LAYER M4 ;
		RECT 155.983 121.019 159.941 121.071 ;
		LAYER M4 ;
		RECT 155.983 121.253 159.941 121.305 ;
		LAYER M4 ;
		RECT 155.983 125.051 159.941 125.103 ;
		LAYER M4 ;
		RECT 155.983 125.285 159.941 125.337 ;
		LAYER M4 ;
		RECT 155.983 129.083 159.941 129.135 ;
		LAYER M4 ;
		RECT 155.983 129.317 159.941 129.369 ;
		LAYER M4 ;
		RECT 155.983 133.115 159.941 133.167 ;
		LAYER M4 ;
		RECT 155.983 133.349 159.941 133.401 ;
		LAYER M4 ;
		RECT 155.983 137.147 159.941 137.199 ;
		LAYER M4 ;
		RECT 155.983 137.381 159.941 137.433 ;
		LAYER M4 ;
		RECT 155.983 141.179 159.941 141.231 ;
		LAYER M4 ;
		RECT 155.983 141.413 159.941 141.465 ;
		LAYER M4 ;
		RECT 208.268 57.539 211.373 57.589 ;
		LAYER M4 ;
		RECT 208.268 58.767 209.663 58.817 ;
		LAYER M4 ;
		RECT 210.555 61.531 211.366 61.629 ;
		LAYER M4 ;
		RECT 210.555 69.087 218.835 69.185 ;
		LAYER M4 ;
		RECT 214.699 73.557 217.574 73.655 ;
		LAYER M4 ;
		RECT 217.492 71.858 218.736 71.908 ;
		LAYER M4 ;
		RECT 218.686 71.725 218.835 71.775 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 220.677 144.672 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 220.677 144.672 ;
	END
END TS1N16FFCLLSVTA8192X32M8SW

END LIBRARY
