**** Created by MC2: Version 2013.12.00.f on 2025/06/23, 08:27:51 

************************************************************************
* auCdl Netlist:
* 
* Library Name:  N16_FFC_CHAR_MB_BOS
* Top Cell Name: LEAFCELLS
* View Name:     schematic
* Netlisted on:  Jan  5 14:07:37 2017
************************************************************************

*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.PARAM


*.PIN vss
.SUBCKT ndio_mac PLUS MINUS 
.ENDS

************************************************************************
* Library Name: TSMC  
* Cell Name:    nand2_svt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC    
* Cell Name:    nand2_ulvt_mac_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_nand2_ulvt_mac_pcell_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
MM2 TSMC_7 TSMC_2 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_7 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_8 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_8 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: tsmcN16
* Cell Name:    inv_lvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_inv_lvt_mac_pcell_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_4:O 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_lvt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_lvt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC  
* Cell Name:    inv_svt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_4:O 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC    
* Cell Name:    inv_ulvt_macN_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_4:O 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC    
* Cell Name:    inv_ulvt_mac_pcell_1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_4:O 
MM1 TSMC_4 TSMC_3 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_4 TSMC_3 TSMC_1 TSMC_2 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC  
* Cell Name:    nand3_svt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_nand3_svt_mac_pcell_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I 
*.PININFO  TSMC_8:O 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC    
* Cell Name:    nand3_ulvt_mac_pcell_2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_nand3_ulvt_mac_pcell_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I 
*.PININFO  TSMC_8:O 
MM3 TSMC_8 TSMC_3 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_8 TSMC_2 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_6 TSMC_7 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM6 TSMC_9 TSMC_3 TSMC_4 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_10 TSMC_2 TSMC_9 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_10 TSMC_5 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    PRECHARGE_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_PRECHARGE_M8 TSMC_1 TSMC_2 TSMC_3 VDDAI VDDI 
*.PININFO  TSMC_3:I TSMC_1:B TSMC_2:B VDDAI:B VDDI:B 
MP0_MIXV_USD VDDAI TSMC_3 TSMC_1 VDDI pch_svt_mac l=20n nfin=8 m=1 
MP5_MIXV_USD TSMC_1 TSMC_3 TSMC_2 VDDI pch_svt_mac l=20n nfin=3 m=1 
MP17_MIXV_USD TSMC_2 TSMC_3 VDDAI VDDI pch_svt_mac l=20n nfin=8 m=1 
.ENDS

************************************************************************
* Library Name: TSMC  
* Cell Name:    nor2_svt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_svt_mac l=p_l nfin=p_nfin m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_svt_mac l=n_l nfin=n_nfin m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC    
* Cell Name:    nor2_ulvt_mac_pcell_3
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_nor2_ulvt_mac_pcell_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
MM2 TSMC_7 TSMC_2 TSMC_8 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_8 TSMC_1 TSMC_5 TSMC_6 pch_ulvt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_7 TSMC_2 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_7 TSMC_1 TSMC_3 TSMC_4 nch_ulvt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    TKBL_TRKPRE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_TKBL_TRKPRE TSMC_1 TSMC_2 TSMC_3 VDDAI VDDI VSSI 
+ TSMC_4 TSMC_5 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_4:O TSMC_5:O TSMC_2:B VDDAI:B VDDI:B VSSI:B 
MM02 TSMC_5 TSMC_6 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MM01 TSMC_5 TSMC_6 VSSI VSSI nch_svt_mac l=20n nfin=12 m=1 
MM2 TSMC_7 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_7 TSMC_6 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MM1 TSMC_3 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_4 TSMC_7 VDDAI VDDI pch_svt_mac l=20n nfin=17 m=2 
MM8 TSMC_6 TSMC_6 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_2 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=6 m=2 
MM4 TSMC_6 TSMC_7 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: TSMC  
* Cell Name:    nor3_svt_mac_pcell_4
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_nor3_svt_mac_pcell_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I 
*.PININFO  TSMC_8:O 
MM3 TSMC_8 TSMC_3 TSMC_9 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM2 TSMC_9 TSMC_2 TSMC_10 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_10 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM6 TSMC_8 TSMC_3 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM5 TSMC_8 TSMC_2 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM4 TSMC_8 TSMC_1 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: TSMC  
* Cell Name:    tri_svt_mac_pcell_5
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I 
*.PININFO  TSMC_8:O 
MM2 TSMC_8 TSMC_3 TSMC_9 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM1 TSMC_9 TSMC_1 TSMC_6 TSMC_7 pch_svt_mac l=p_l nfin=p_nfin 
+ m=p_totalM 
MM4 TSMC_10 TSMC_1 TSMC_4 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
MM3 TSMC_8 TSMC_2 TSMC_10 TSMC_5 nch_svt_mac l=n_l nfin=n_nfin 
+ m=n_totalM 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_WLP_S_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_WLP_S_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 VDDAI VDDHD VDDI VSSI TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 TSMC_14 
*.PININFO  TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_8:I 
*.PININFO  TSMC_9:I TSMC_14:I TSMC_1:O TSMC_2:O TSMC_10:O TSMC_11:O TSMC_12:O 
*.PININFO  TSMC_13:O VDDAI:B VDDHD:B VDDI:B VSSI:B 
MM35 TSMC_15 TSMC_7 TSMC_16 VSSI nch_svt_mac l=16.0n nfin=10 m=4 
MM34 TSMC_17 TSMC_6 TSMC_16 VSSI nch_svt_mac l=16.0n nfin=10 m=4 
MM32 TSMC_18 TSMC_5 TSMC_16 VSSI nch_svt_mac l=16.0n nfin=10 m=4 
MM28 TSMC_19 TSMC_4 TSMC_16 VSSI nch_svt_mac l=16.0n nfin=10 m=4 
MM36 TSMC_20 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN0_MIXV_ULVT TSMC_20 TSMC_21 TSMC_22 VSSI nch_ulvt_mac l=16.0n nfin=9 
+ m=3 
MN1_MIXV_ULVT TSMC_22 TSMC_23 VSSI VSSI nch_ulvt_mac l=16.0n nfin=9 m=3 
MM2 TSMC_1 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM0_MIXV_ULVT TSMC_16 TSMC_3 VSSI VSSI nch_ulvt_mac l=16.0n nfin=7 m=10 
MP0_MIXV_ULVT TSMC_20 TSMC_21 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=10 
+ m=3 
MP1 TSMC_20 TSMC_23 VDDHD VDDI pch_svt_mac l=16.0n nfin=6 m=1 
MM16_MIXV_ULVT TSMC_17 TSMC_3 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 
+ m=3 
MM9_MIXV_ULVT TSMC_18 TSMC_3 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 m=3 
MM20_MIXV_ULVT TSMC_19 TSMC_3 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 
+ m=3 
MM15_MIXV_ULVT TSMC_15 TSMC_7 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 
+ m=1 
MM13_MIXV_ULVT TSMC_17 TSMC_6 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 
+ m=1 
MM12_MIXV_ULVT TSMC_19 TSMC_4 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 
+ m=1 
MM10_MIXV_ULVT TSMC_18 TSMC_5 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 
+ m=1 
MM21_MIXV_ULVT TSMC_15 TSMC_3 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=6 
+ m=3 
XI543_MIXV_ULVT_N VSSI VSSI TSMC_20 TSMC_1 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=8 n_nfin=11 n_l=16.0n 
+ p_totalM=12 p_nfin=12 p_l=16.0n 
XI550 VSSI VSSI TSMC_24 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI571_MIXV_ULVT VSSI VSSI TSMC_3 TSMC_21 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=2 n_nfin=5 n_l=16.0n 
+ p_totalM=1 p_nfin=4 p_l=16.0n 
XI532_MIXV_ULVT_N VSSI VSSI TSMC_18 TSMC_11 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=10 n_nfin=7 n_l=16.0n 
+ p_totalM=10 p_nfin=11 p_l=16.0n 
XI531_MIXV_ULVT_N VSSI VSSI TSMC_15 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=10 n_nfin=7 n_l=16.0n 
+ p_totalM=10 p_nfin=11 p_l=16.0n 
XI533_MIXV_ULVT_N VSSI VSSI TSMC_17 TSMC_12 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=10 n_nfin=7 n_l=16.0n 
+ p_totalM=10 p_nfin=11 p_l=16.0n 
XI534_MIXV_ULVT_N VSSI VSSI TSMC_19 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=10 n_nfin=7 n_l=16.0n 
+ p_totalM=10 p_nfin=11 p_l=16.0n 
XI551 TSMC_20 TSMC_20 TSMC_20 VSSI VSSI VDDHD VDDI TSMC_24 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI577 TSMC_21 TSMC_21 TSMC_21 VSSI VSSI VDDHD VDDI TSMC_25 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI570 TSMC_25 TSMC_25 TSMC_25 VSSI VSSI VDDHD VDDI TSMC_23 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_Y4_LG_M16
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_Y4_LG_M16 TSMC_1 VDDHD VDDI VSSI TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
*.PININFO  TSMC_8:O TSMC_9:O TSMC_10:O VDDHD:B VDDI:B VSSI:B 
MN3<3> TSMC_10 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN3<2> TSMC_9 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN3<1> TSMC_8 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN3<0> TSMC_7 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN21 TSMC_11 TSMC_2 VSSI VSSI nch_svt_mac l=20n nfin=12 m=1 
MP31 TSMC_11 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM17<3> TSMC_12 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM17<2> TSMC_13 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM17<1> TSMC_14 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM17<0> TSMC_15 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
XI407<3> VSSI VSSI TSMC_12 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=6 n_nfin=10 n_l=20n p_totalM=6 
+ p_nfin=10 p_l=20n 
XI407<2> VSSI VSSI TSMC_13 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=6 n_nfin=10 n_l=20n p_totalM=6 
+ p_nfin=10 p_l=20n 
XI407<1> VSSI VSSI TSMC_14 TSMC_9 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=6 n_nfin=10 n_l=20n p_totalM=6 
+ p_nfin=10 p_l=20n 
XI407<0> VSSI VSSI TSMC_15 TSMC_10 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=6 n_nfin=10 n_l=20n p_totalM=6 
+ p_nfin=10 p_l=20n 
XNA2<3> TSMC_11 VSSI TSMC_3 TSMC_12 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XNA2<2> TSMC_11 VSSI TSMC_4 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XNA2<1> TSMC_11 VSSI TSMC_5 TSMC_14 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XNA2<0> TSMC_11 VSSI TSMC_6 TSMC_15 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=4 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_Y10_NAND3
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_Y10_NAND3 TSMC_1 VDDHD VDDI VSSI TSMC_2 TSMC_3 
+ TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:O 
*.PININFO  TSMC_8:O VDDHD:B VDDI:B VSSI:B 
MM19 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM11 TSMC_10 TSMC_6 VSSI VSSI nch_svt_mac l=20n nfin=10 m=3 
MM13 TSMC_8 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM21 TSMC_11 TSMC_2 TSMC_10 VSSI nch_svt_mac l=20n nfin=10 m=3 
MM15 TSMC_11 TSMC_3 TSMC_10 VSSI nch_svt_mac l=20n nfin=10 m=3 
MM2 TSMC_12 TSMC_4 TSMC_11 VSSI nch_svt_mac l=20n nfin=11 m=1 
MN3 TSMC_7 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_7 TSMC_12 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MM14 TSMC_9 TSMC_5 TSMC_11 VSSI nch_svt_mac l=20n nfin=11 m=1 
MM23 TSMC_13 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM22 TSMC_14 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM20 TSMC_8 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=10 m=10 
MM18 TSMC_9 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM16 TSMC_9 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM3 TSMC_12 TSMC_3 TSMC_13 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM17 TSMC_9 TSMC_3 TSMC_14 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM12 TSMC_12 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM8 TSMC_12 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM4 TSMC_7 TSMC_12 VDDHD VDDI pch_svt_mac l=20n nfin=10 m=10 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_Y10_NAND2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_Y10_NAND2 TSMC_1 VDDHD VDDI VSSI TSMC_2 TSMC_3 
+ TSMC_4 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:O VDDHD:B VDDI:B VSSI:B 
MM11_MIXV_ULVT TSMC_5 TSMC_2 VSSI VSSI nch_ulvt_mac l=16.0n nfin=11 m=1 
MM2_MIXV_ULVT TSMC_6 TSMC_3 TSMC_5 VSSI nch_ulvt_mac l=16.0n nfin=11 m=1 
MN3 TSMC_4 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_4 TSMC_6 VSSI VSSI nch_svt_mac l=20n nfin=10 m=5 
MM3_MIXV_ULVT TSMC_6 TSMC_2 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=4 m=1 
MM8_MIXV_ULVT TSMC_6 TSMC_3 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=4 m=1 
MM4 TSMC_4 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=10 m=6 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_READ_NOR
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_READ_NOR TSMC_1 TSMC_2 TSMC_3 VDDHD VDDI VSSI 
+ TSMC_4 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_3:O VDDHD:B VDDI:B VSSI:B 
MN1 TSMC_5 TSMC_2 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
XI428 VSSI VSSI TSMC_1 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI426 VSSI VSSI TSMC_5 TSMC_3 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=6 n_nfin=10 n_l=20n p_totalM=6 
+ p_nfin=10 p_l=20n 
XI631_MIXV_ULVT TSMC_4 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_5 
+ S1ALLSVTSW2000X20_nor2_ulvt_mac_pcell_3 n_totalM=1 n_nfin=8 n_l=16.0n 
+ p_totalM=1 p_nfin=8 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_Y10
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_Y10 TSMC_1 VDDHD VDDI VSSI TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:O TSMC_6:O VDDHD:B VDDI:B 
*.PININFO  VSSI:B 
MN21 TSMC_7 TSMC_2 VSSI VSSI nch_svt_mac l=20n nfin=8 m=1 
MM2 TSMC_8 TSMC_3 TSMC_7 VSSI nch_svt_mac l=20n nfin=10 m=1 
MM0 TSMC_6 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN3 TSMC_5 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_6 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=10 m=6 
MM5 TSMC_5 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=10 m=6 
MM10 TSMC_9 TSMC_4 TSMC_7 VSSI nch_svt_mac l=20n nfin=10 m=1 
MM9 TSMC_9 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MP31 TSMC_7 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_8 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM6 TSMC_6 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=10 m=6 
MM11 TSMC_9 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM8 TSMC_8 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM4 TSMC_5 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=10 m=6 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    LCTRL_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_LCTRL_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 VDDHD VDDI VSSI 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I 
*.PININFO  TSMC_7:I TSMC_8:I TSMC_9:I TSMC_10:I TSMC_11:I TSMC_12:I 
*.PININFO  TSMC_29:I TSMC_30:I TSMC_33:I TSMC_36:I TSMC_37:I TSMC_38:I 
*.PININFO  TSMC_13:O 
*.PININFO  TSMC_14:O TSMC_15:O TSMC_16:O TSMC_17:O 
*.PININFO  TSMC_18:O TSMC_19:O TSMC_20:O TSMC_21:O 
*.PININFO  TSMC_22:O TSMC_23:O TSMC_24:O TSMC_25:O 
*.PININFO  TSMC_26:O TSMC_27:O TSMC_28:O TSMC_31:O TSMC_32:O 
*.PININFO  TSMC_34:O TSMC_35:O TSMC_39:O TSMC_40:O VDDHD:B VDDI:B VSSI:B 
XNOR0_MIXV_ULVT TSMC_4 TSMC_3 VSSI VSSI VDDHD VDDI TSMC_41 
+ S1ALLSVTSW2000X20_nor2_ulvt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XXDRV_Y4_D<0> TSMC_29 VDDHD VDDI VSSI TSMC_42 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ S1ALLSVTSW2000X20_XDRV_Y4_LG_M16 
XXDRV_Y4_D<1> TSMC_29 VDDHD VDDI VSSI TSMC_42 TSMC_9 TSMC_10 TSMC_11 
+ TSMC_12 TSMC_17 TSMC_18 TSMC_19 TSMC_20 
+ S1ALLSVTSW2000X20_XDRV_Y4_LG_M16 
XXDRV_Y4_U<0> TSMC_29 VDDHD VDDI VSSI TSMC_43 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ S1ALLSVTSW2000X20_XDRV_Y4_LG_M16 
XXDRV_Y4_U<1> TSMC_29 VDDHD VDDI VSSI TSMC_43 TSMC_9 TSMC_10 TSMC_11 
+ TSMC_12 TSMC_25 TSMC_26 TSMC_27 TSMC_28 
+ S1ALLSVTSW2000X20_XDRV_Y4_LG_M16 
XXDRV_W TSMC_29 VDDHD VDDI VSSI TSMC_3 TSMC_4 TSMC_37 TSMC_38 TSMC_33 
+ TSMC_34 TSMC_35 S1ALLSVTSW2000X20_XDRV_Y10_NAND3 
XXDRV_R TSMC_29 VDDHD VDDI VSSI TSMC_44 TSMC_30 TSMC_31 
+ S1ALLSVTSW2000X20_XDRV_Y10_NAND2 
XXDRV_READ TSMC_44 TSMC_29 TSMC_32 VDDHD VDDI VSSI TSMC_36 
+ S1ALLSVTSW2000X20_XDRV_READ_NOR 
XXDRV_YL TSMC_29 VDDHD VDDI VSSI TSMC_44 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ S1ALLSVTSW2000X20_XDRV_Y10 
XD3_BUF_MIXV_ULVT<1> VSSI VSSI TSMC_4 TSMC_45 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=1 n_nfin=5 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XD3_BUF_MIXV_ULVT<0> VSSI VSSI TSMC_3 TSMC_46 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=1 n_nfin=5 n_l=16.0n 
+ p_totalM=1 p_nfin=3 p_l=16.0n 
XI252_MIXV_ULVT<1> VSSI VSSI TSMC_45 TSMC_43 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=2 n_nfin=3 n_l=16.0n 
+ p_totalM=2 p_nfin=8 p_l=16.0n 
XI252_MIXV_ULVT<0> VSSI VSSI TSMC_46 TSMC_42 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=2 n_nfin=3 n_l=16.0n 
+ p_totalM=2 p_nfin=8 p_l=16.0n 
XINV4 VSSI VSSI TSMC_47 TSMC_48 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV5 VSSI VSSI TSMC_48 TSMC_49 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV0 VSSI VSSI TSMC_41 TSMC_50 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV3 VSSI VSSI TSMC_51 TSMC_47 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV2 VSSI VSSI TSMC_52 TSMC_51 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV1 VSSI VSSI TSMC_50 TSMC_52 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XNAND0_MIXV_ULVT TSMC_52 TSMC_41 VSSI VSSI VDDHD VDDI TSMC_44 
+ S1ALLSVTSW2000X20_nand2_ulvt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=16.0n 
+ p_totalM=1 p_nfin=8 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    SA_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_SA_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDDAI VDDI VSSI 
*.PININFO  TSMC_7:I TSMC_8:I TSMC_9:I TSMC_10:I TSMC_1:B TSMC_2:B TSMC_3:B 
*.PININFO  TSMC_4:B 
*.PININFO  TSMC_5:B TSMC_6:B VDDAI:B VDDI:B VSSI:B 
MN0_MIXV_USD TSMC_11 TSMC_12 TSMC_13 VSSI nch_svt_mac l=20n nfin=10 m=4 
MN1_MIXV_USD TSMC_12 TSMC_11 TSMC_13 VSSI nch_svt_mac l=20n nfin=10 m=4 
MN11 TSMC_5 TSMC_14 VSSI VSSI nch_svt_mac l=20n nfin=10 m=3 
MM0 TSMC_6 TSMC_15 VSSI VSSI nch_svt_mac l=20n nfin=10 m=3 
MN2_MIXV_USD TSMC_13 TSMC_10 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MP2_MIXV_SULVT TSMC_11 TSMC_12 VDDAI VDDI pch_ulvt_mac l=20n nfin=5 m=1 
MP6_MIXV_SULVT TSMC_4 TSMC_8 TSMC_11 VDDI pch_ulvt_mac l=20n nfin=5 m=1 
MP7_MIXV_SULVT TSMC_2 TSMC_8 TSMC_12 VDDI pch_ulvt_mac l=20n nfin=5 m=1 
MP13_MIXV_SULVT TSMC_3 TSMC_7 TSMC_11 VDDI pch_ulvt_mac l=20n nfin=5 
+ m=1 
MP14_MIXV_SULVT TSMC_1 TSMC_7 TSMC_12 VDDI pch_ulvt_mac l=20n nfin=5 
+ m=1 
MP3_MIXV_SULVT TSMC_12 TSMC_11 VDDAI VDDI pch_ulvt_mac l=20n nfin=5 m=1 
MP8_MIXV_SULVT TSMC_11 TSMC_9 TSMC_12 VDDI pch_ulvt_mac l=20n nfin=5 
+ m=2 
MP11_MIXV_SULVT TSMC_12 TSMC_9 VDDAI VDDI pch_ulvt_mac l=20n nfin=5 m=1 
MP10_MIXV_SULVT TSMC_11 TSMC_9 VDDAI VDDI pch_ulvt_mac l=20n nfin=5 m=1 
XINV1 VSSI VSSI TSMC_12 TSMC_15 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XINV0 VSSI VSSI TSMC_11 TSMC_14 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    IO_RWBLK_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_IO_RWBLK_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 VDDAI 
+ VDDI VSSI TSMC_16 TSMC_17 TSMC_18 TSMC_19 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_11:I TSMC_12:I TSMC_13:I 
*.PININFO  TSMC_15:I 
*.PININFO  TSMC_17:I TSMC_14:O TSMC_16:O TSMC_18:O TSMC_19:O TSMC_5:B TSMC_6:B 
*.PININFO  TSMC_7:B TSMC_8:B 
*.PININFO  TSMC_9:B TSMC_10:B VDDAI:B VDDI:B VSSI:B 
XSA TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ VDDAI VDDI VSSI S1ALLSVTSW2000X20_SA_M8 
MN0_MIXV_UWAS TSMC_16 TSMC_11 VSSI VSSI nch_ulvt_mac l=20n nfin=10 m=4 
MN13_MIXV_UWAS TSMC_19 TSMC_12 VSSI VSSI nch_ulvt_mac l=20n nfin=10 m=4 
MM3_MIXV_DFTUUU TSMC_24 TSMC_25 VSSI VSSI nch_ulvt_mac l=20n nfin=4 m=1 
XI49 TSMC_26 TSMC_25 VSSI VSSI VDDAI VDDI TSMC_22 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n 
+ p_totalM=1 p_nfin=3 p_l=20n 
MP25 TSMC_19 TSMC_12 VDDAI VDDI pch_svt_mac l=20n nfin=7 m=1 
MP27 TSMC_16 TSMC_11 VDDAI VDDI pch_svt_mac l=20n nfin=7 m=1 
MM1 TSMC_21 TSMC_25 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MM2 TSMC_20 TSMC_25 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
XINV5 VSSI VSSI TSMC_26 TSMC_27 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=3 p_l=20n 
XI47_MIXV_ULVT_N VSSI VSSI TSMC_13 TSMC_26 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=1 n_nfin=4 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
XI273_MIXV_ULVT_N TSMC_24 VSSI TSMC_1 TSMC_20 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=1 n_nfin=4 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
XI108 VSSI VSSI TSMC_23 TSMC_25 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI1 VSSI VSSI TSMC_17 TSMC_28 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI111 VSSI VSSI TSMC_26 TSMC_14 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI268 VSSI VSSI TSMC_28 TSMC_18 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI248 VSSI VSSI TSMC_15 TSMC_23 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI272_MIXV_ULVT_N TSMC_24 VSSI TSMC_2 TSMC_21 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_macN_pcell_1 n_totalM=1 n_nfin=4 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DOUT_INV
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DOUT_INV TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDDHD VDDI VSSI TSMC_7 TSMC_8 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_6:I TSMC_7:I TSMC_8:I TSMC_5:O TSMC_3:B 
*.PININFO  TSMC_4:B 
*.PININFO  VDDHD:B VDDI:B VSSI:B 
MP7_MIXV_ULVT TSMC_4 TSMC_9 VDDHD VDDI pch_ulvt_mac l=20n nfin=10 m=3 
MP6_MIXV_ULVT TSMC_3 TSMC_4 VDDHD VDDI pch_ulvt_mac l=20n nfin=2 m=1 
MM3_MIXV_ULVT TSMC_10 TSMC_6 VDDHD VDDI pch_ulvt_mac l=20n nfin=6 m=4 
MM2_MIXV_ULVT TSMC_5 TSMC_11 TSMC_10 VDDI pch_ulvt_mac l=20n nfin=6 m=4 
MP8_MIXV_ULVT TSMC_3 TSMC_9 VDDHD VDDI pch_ulvt_mac l=20n nfin=10 m=3 
MP0_MIXV_ULVT TSMC_4 TSMC_3 VDDHD VDDI pch_ulvt_mac l=20n nfin=2 m=1 
MM41_MIXV_ULVT TSMC_12 TSMC_9 VSSI VSSI nch_ulvt_mac l=20n nfin=6 m=1 
MM40_MIXV_ULVT TSMC_3 TSMC_13 TSMC_12 VSSI nch_ulvt_mac l=16.0n nfin=5 
+ m=1 
MM39_MIXV_ULVT TSMC_2 TSMC_6 VSSI VSSI nch_ulvt_mac l=20n nfin=2 m=1 
MM33_MIXV_ULVT TSMC_5 TSMC_6 VSSI VSSI nch_ulvt_mac l=20n nfin=2 m=1 
MM0_MIXV_ULVT TSMC_5 TSMC_11 VSSI VSSI nch_ulvt_mac l=20n nfin=8 m=2 
MM42_MIXV_ULVT TSMC_4 TSMC_14 TSMC_12 VSSI nch_ulvt_mac l=16.0n nfin=5 
+ m=1 
XI180_MIXV_ULVT TSMC_15 TSMC_3 VSSI VSSI VDDHD VDDI TSMC_11 
+ S1ALLSVTSW2000X20_nand2_ulvt_mac_pcell_0 n_totalM=1 n_nfin=5 n_l=16.0n 
+ p_totalM=1 p_nfin=5 p_l=16.0n 
XI181_MIXV_ULVT TSMC_4 TSMC_11 VSSI VSSI VDDHD VDDI TSMC_15 
+ S1ALLSVTSW2000X20_nand2_ulvt_mac_pcell_0 n_totalM=1 n_nfin=5 n_l=16.0n 
+ p_totalM=1 p_nfin=2 p_l=16.0n 
XI166 VSSI VSSI TSMC_2 TSMC_16 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI168_MIXV_ULVT VSSI VSSI TSMC_3 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI169_MIXV_ULVT VSSI VSSI TSMC_4 TSMC_14 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI176 VSSI VSSI TSMC_7 TSMC_17 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI95 TSMC_1 TSMC_6 VSSI VSSI VDDI VDDI TSMC_18 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI160 TSMC_17 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_9 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=9 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DIN_NM
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DIN_NM TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VDDHD VDDI VSSI 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_4:I TSMC_7:I TSMC_1:O TSMC_5:O TSMC_6:O 
*.PININFO  VDDHD:B VDDI:B VSSI:B 
MM29 TSMC_8 TSMC_9 TSMC_10 VDDI pch_svt_mac l=20n nfin=2 m=1 
MP10 TSMC_11 TSMC_12 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MM51 TSMC_13 TSMC_14 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MM52 TSMC_11 TSMC_15 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MM28 TSMC_10 TSMC_15 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM26 TSMC_16 TSMC_12 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM53 TSMC_11 TSMC_17 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MM39 TSMC_18 TSMC_17 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM27 TSMC_8 TSMC_19 TSMC_16 VDDI pch_svt_mac l=20n nfin=2 m=1 
MP2 TSMC_1 TSMC_20 TSMC_21 VDDI pch_svt_mac l=20n nfin=2 m=1 
MP1 TSMC_13 TSMC_12 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP5 TSMC_1 TSMC_4 TSMC_22 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM40 TSMC_23 TSMC_9 TSMC_18 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM38 TSMC_24 TSMC_12 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM41 TSMC_23 TSMC_25 TSMC_24 VDDI pch_svt_mac l=20n nfin=2 m=1 
MP4 TSMC_22 TSMC_26 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM54 TSMC_13 TSMC_17 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP3 TSMC_21 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM45 TSMC_23 TSMC_12 TSMC_27 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM35 TSMC_8 TSMC_12 TSMC_28 VSSI nch_svt_mac l=20n nfin=2 m=1 
MN1 TSMC_11 TSMC_15 TSMC_29 VSSI nch_svt_mac l=20n nfin=3 m=2 
MM44 TSMC_27 TSMC_17 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM42 TSMC_23 TSMC_25 TSMC_30 VSSI nch_svt_mac l=20n nfin=2 m=1 
MN33 TSMC_13 TSMC_14 TSMC_29 VSSI nch_svt_mac l=20n nfin=6 m=1 
MM37 TSMC_28 TSMC_15 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM43 TSMC_30 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN13 TSMC_31 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM34 TSMC_8 TSMC_19 TSMC_32 VSSI nch_svt_mac l=20n nfin=2 m=1 
MN4 TSMC_31 TSMC_26 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN6 TSMC_1 TSMC_20 TSMC_31 VSSI nch_svt_mac l=20n nfin=2 m=1 
MN2 TSMC_29 TSMC_12 TSMC_33 VSSI nch_svt_mac l=20n nfin=5 m=2 
MM36 TSMC_32 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MN7 TSMC_33 TSMC_17 VSSI VSSI nch_svt_mac l=20n nfin=10 m=4 
MN5 TSMC_1 TSMC_2 TSMC_31 VSSI nch_svt_mac l=20n nfin=2 m=1 
XI339 TSMC_7 TSMC_23 VSSI VSSI VDDHD VDDI TSMC_17 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI329 VSSI VSSI TSMC_8 TSMC_15 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI317_MIXV_DFTUUU VSSI VSSI TSMC_9 TSMC_12 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI357 VSSI VSSI TSMC_34 TSMC_19 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI358 VSSI VSSI TSMC_35 TSMC_25 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI367 VSSI VSSI TSMC_2 TSMC_35 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI331 VSSI VSSI TSMC_15 TSMC_14 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI325 VSSI VSSI TSMC_2 TSMC_26 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI314_MIXV_DFTUUU VSSI VSSI TSMC_3 TSMC_9 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI366 VSSI VSSI TSMC_4 TSMC_34 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI332 VSSI VSSI TSMC_11 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=5 n_nfin=4 n_l=20n p_totalM=4 
+ p_nfin=10 p_l=20n 
XI333 VSSI VSSI TSMC_13 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=5 n_nfin=4 n_l=20n p_totalM=5 
+ p_nfin=8 p_l=20n 
XI321 VSSI VSSI TSMC_4 TSMC_20 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    IO_INV_NM
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_IO_INV_NM TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 VDDHD VDDI VSSI TSMC_11 TSMC_12 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_10:I TSMC_11:I TSMC_12:I 
*.PININFO  TSMC_7:O TSMC_8:O 
*.PININFO  TSMC_9:O TSMC_5:B TSMC_6:B VDDHD:B VDDI:B VSSI:B 
XDOUT TSMC_1 TSMC_13 TSMC_5 TSMC_6 TSMC_9 TSMC_10 VDDHD VDDI VSSI TSMC_11 
+ TSMC_12 S1ALLSVTSW2000X20_DOUT_INV 
XDIN TSMC_13 TSMC_2 TSMC_3 TSMC_4 TSMC_7 TSMC_8 TSMC_10 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DIN_NM 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    TM_BUF
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_TM_BUF TSMC_1 TSMC_2 TSMC_3 VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_3:I VDDHD:I VDDI:I VSSI:I TSMC_2:O 
XINV0 VSSI VSSI TSMC_1 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI12 TSMC_4 TSMC_3 VSSI VSSI VDDI VDDI TSMC_2 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    RWA_TSEL
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_RWA_TSEL TSMC_1 TSMC_2 TSMC_3 VDDHD VDDI VSSI TSMC_4 
+ TSMC_5 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:O TSMC_5:O VDDHD:B VDDI:B VSSI:B 
MM11 TSMC_6 TSMC_7 TSMC_8 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM8 TSMC_8 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_7 TSMC_9 TSMC_10 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_10 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_11 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM0 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM10 TSMC_6 TSMC_7 TSMC_12 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM9 TSMC_12 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM6 TSMC_7 TSMC_9 TSMC_13 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_13 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_9 TSMC_1 TSMC_14 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM2 TSMC_14 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
XI2 TSMC_1 TSMC_5 VSSI VSSI VDDHD VDDI TSMC_15 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI1 TSMC_15 TSMC_16 VSSI VSSI VDDHD VDDI TSMC_4 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI0 TSMC_6 TSMC_17 VSSI VSSI VDDHD VDDI TSMC_5 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI4 VSSI VSSI TSMC_2 TSMC_16 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI3 VSSI VSSI TSMC_3 TSMC_17 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    MCTRL_RWA_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_MCTRL_RWA_M8 TSMC_1 TSMC_2 TSMC_3 VDDHD VDDI VSSI 
+ TSMC_4 TSMC_5 TSMC_6 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_1:O VDDHD:B 
*.PININFO  VDDI:B VSSI:B 
XI0 TSMC_3 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_7 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
XI2 TSMC_8 TSMC_9 TSMC_7 VSSI VSSI VDDHD VDDI TSMC_10 
+ S1ALLSVTSW2000X20_nor3_svt_mac_pcell_4 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI3 VSSI VSSI TSMC_10 TSMC_1 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=4 n_nfin=3 n_l=20n p_totalM=4 
+ p_nfin=3 p_l=20n 
MM0 TSMC_10 TSMC_2 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
XI1 TSMC_7 TSMC_4 TSMC_5 VDDHD VDDI VSSI TSMC_8 TSMC_9 
+ S1ALLSVTSW2000X20_RWA_TSEL 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    VHILO
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_VHILO VDDI TSMC_1 TSMC_2 VSSI 
*.PININFO  TSMC_1:O TSMC_2:O VDDI:B VSSI:B 
MN3 VSSI TSMC_3 TSMC_4 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN0 VSSI TSMC_4 TSMC_4 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1 VSSI TSMC_3 TSMC_2 VSSI nch_svt_mac l=20n nfin=9 m=4 
MP7 TSMC_3 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP2 TSMC_1 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=9 m=4 
MP0 TSMC_3 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    PMCTRL_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_PMCTRL_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_2:O TSMC_4:O TSMC_7:O 
*.PININFO  VDDI:B 
*.PININFO  VSSI:B 
XI74 TSMC_8 TSMC_9 VSSI VSSI VDDI VDDI TSMC_10 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI95 TSMC_11 TSMC_5 VSSI VSSI VDDI VDDI TSMC_12 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI97 TSMC_8 TSMC_1 VSSI VSSI VDDI VDDI TSMC_9 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI76 TSMC_6 TSMC_10 TSMC_8 VSSI VSSI VDDI VDDI TSMC_13 
+ S1ALLSVTSW2000X20_nor3_svt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI87 VSSI VSSI TSMC_12 TSMC_7 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=4 n_nfin=10 n_l=20n p_totalM=4 
+ p_nfin=4 p_l=20n 
XI85 VSSI VSSI TSMC_14 TSMC_2 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=4 n_nfin=4 n_l=20n p_totalM=4 
+ p_nfin=8 p_l=20n 
XI86 VSSI VSSI TSMC_13 TSMC_11 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI93 VSSI VSSI TSMC_10 TSMC_14 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI48 VSSI VSSI TSMC_3 TSMC_15 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI94 VSSI VSSI TSMC_8 TSMC_16 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI49 VSSI VSSI TSMC_15 TSMC_8 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=8 p_l=20n 
XI80 VSSI VSSI TSMC_16 TSMC_4 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=4 n_nfin=4 n_l=20n p_totalM=4 
+ p_nfin=8 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    CKG
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_CKG TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ VDDHD VDDI VSSI 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_1:O TSMC_4:O 
*.PININFO  VDDHD:B VDDI:B VSSI:B 
XINV0 TSMC_8 TSMC_6 VSSI VSSI VDDI VDDI TSMC_4 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
XNAND0 TSMC_2 TSMC_7 VSSI VSSI VDDHD VDDI TSMC_9 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n 
+ p_totalM=1 p_nfin=3 p_l=20n 
XNAND3 TSMC_10 TSMC_11 VSSI VSSI VDDHD VDDI TSMC_8 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n 
+ p_totalM=1 p_nfin=3 p_l=20n 
XNAND5 TSMC_4 TSMC_1 VSSI VSSI VDDHD VDDI TSMC_12 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=20n 
+ p_totalM=1 p_nfin=4 p_l=20n 
XNAND2 TSMC_2 TSMC_8 VSSI VSSI VDDHD VDDI TSMC_10 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=3 n_l=20n 
+ p_totalM=1 p_nfin=3 p_l=20n 
XNAND4 TSMC_12 TSMC_13 VSSI VSSI VDDHD VDDI TSMC_1 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=2 n_nfin=5 n_l=20n 
+ p_totalM=2 p_nfin=7 p_l=20n 
XNAND1 TSMC_9 TSMC_1 TSMC_5 VSSI VSSI VDDHD VDDI TSMC_11 
+ S1ALLSVTSW2000X20_nand3_svt_mac_pcell_2 n_totalM=1 n_nfin=3 n_l=20n 
+ p_totalM=1 p_nfin=3 p_l=20n 
XNAND12 TSMC_4 TSMC_3 TSMC_2 VSSI VSSI VDDHD VDDI TSMC_13 
+ S1ALLSVTSW2000X20_nand3_svt_mac_pcell_2 n_totalM=1 n_nfin=7 n_l=20n 
+ p_totalM=1 p_nfin=4 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    RESETD_TSEL_WT_NOR
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_RESETD_TSEL_WT_NOR TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ TSMC_3 TSMC_4 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_4:I TSMC_2:O VDDHD:B VDDI:B VSSI:B 
MM15 TSMC_5 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM14 TSMC_7 TSMC_6 TSMC_5 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM13 TSMC_8 TSMC_9 TSMC_10 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM12 TSMC_10 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM8 TSMC_11 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_12 TSMC_1 TSMC_13 VDDI pch_svt_mac l=20n nfin=5 m=2 
MM0 TSMC_12 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
MM9 TSMC_9 TSMC_1 TSMC_11 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM3 TSMC_13 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
MM17 TSMC_14 TSMC_6 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM16 TSMC_7 TSMC_6 TSMC_14 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM11 TSMC_8 TSMC_9 TSMC_15 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM6 TSMC_12 TSMC_1 TSMC_16 VSSI nch_svt_mac l=20n nfin=5 m=1 
MM2 TSMC_16 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=5 m=1 
MM7 TSMC_9 TSMC_1 TSMC_17 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_17 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_12 TSMC_7 TSMC_16 VSSI nch_svt_mac l=20n nfin=5 m=1 
MM10 TSMC_15 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
XI90 TSMC_8 TSMC_4 VSSI VSSI VDDHD VDDI TSMC_6 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=20n 
+ p_totalM=1 p_nfin=3 p_l=20n 
XI574 TSMC_12 TSMC_6 VSSI VSSI VDDHD VDDI TSMC_2 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=20n 
+ p_totalM=1 p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    RESETD_TSEL_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_RESETD_TSEL_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ VDDHD VDDI VSSI TSMC_6 TSMC_7 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:O TSMC_7:O 
*.PININFO  VDDHD:B VDDI:B 
*.PININFO  VSSI:B 
MM3 TSMC_8 TSMC_9 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM2 TSMC_10 TSMC_9 TSMC_8 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM10 TSMC_11 TSMC_10 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM9 TSMC_12 TSMC_10 TSMC_11 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM22 TSMC_13 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM16 TSMC_9 TSMC_1 TSMC_13 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM8 TSMC_14 TSMC_10 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_12 TSMC_10 TSMC_15 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_16 TSMC_9 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM6 TSMC_15 TSMC_10 TSMC_14 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM0 TSMC_10 TSMC_9 TSMC_17 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_17 TSMC_9 TSMC_16 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_18 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM31 TSMC_19 TSMC_1 TSMC_18 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM30 TSMC_9 TSMC_1 TSMC_19 VDDI pch_svt_mac l=20n nfin=2 m=1 
XND5 TSMC_5 TSMC_12 VSSI VSSI VDDHD VDDI TSMC_7 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
XND1_MIXV_ULVT TSMC_4 TSMC_20 VSSI VSSI VDDHD VDDI TSMC_6 
+ S1ALLSVTSW2000X20_nand2_ulvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=16.0n 
+ p_totalM=1 p_nfin=2 p_l=16.0n 
XND0_MIXV_ULVT TSMC_7 TSMC_21 VSSI VSSI VDDHD VDDI TSMC_20 
+ S1ALLSVTSW2000X20_nand2_ulvt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=16.0n 
+ p_totalM=1 p_nfin=2 p_l=16.0n 
XI79_MIXV_SLL VSSI VSSI TSMC_22 TSMC_21 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_lvt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=16.0n 
+ p_totalM=1 p_nfin=2 p_l=16.0n 
XI599_MIXV_SUL2 VSSI VSSI TSMC_1 TSMC_22 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_lvt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=16.0n 
+ p_totalM=1 p_nfin=2 p_l=16.0n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    RESETD_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_RESETD_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 VDDHD VDDI VSSI TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_6:I TSMC_9:I TSMC_10:I TSMC_11:I TSMC_13:I 
*.PININFO  TSMC_17:I TSMC_18:I 
*.PININFO  TSMC_19:I TSMC_20:I TSMC_21:I TSMC_22:I TSMC_23:I TSMC_1:O TSMC_4:O 
*.PININFO  TSMC_5:O TSMC_7:O TSMC_8:O TSMC_14:O TSMC_16:O TSMC_12:B 
*.PININFO  VDDHD:B VDDI:B VSSI:B TSMC_15:B 
XI635 TSMC_24 TSMC_25 VDDHD VDDI VSSI TSMC_22 TSMC_23 
+ S1ALLSVTSW2000X20_RESETD_TSEL_WT_NOR 
XI630 TSMC_26 TSMC_27 VDDHD VDDI VSSI TSMC_20 TSMC_21 
+ S1ALLSVTSW2000X20_RESETD_TSEL_WT_NOR 
MM19_MIXV_DFTUUU TSMC_28 TSMC_26 VDDHD VDDI pch_ulvt_mac l=16.0n nfin=7 
+ m=2 
MM3_MIXV_WLDV TSMC_1 TSMC_29 VDDHD VDDI pch_svt_mac l=20n nfin=11 m=3 
MM20 TSMC_30 TSMC_31 TSMC_24 VDDI pch_svt_mac l=16.0n nfin=4 m=2 
MP16 TSMC_14 TSMC_32 VDDI VDDI pch_svt_mac l=16.0n nfin=4 m=11 
MM0 TSMC_12 TSMC_33 TSMC_24 VDDI pch_svt_mac l=16.0n nfin=4 m=2 
MM2_MIXV_DFTUUU TSMC_34 TSMC_27 TSMC_28 VDDI pch_ulvt_mac l=16.0n 
+ nfin=7 m=2 
XI636 TSMC_35 TSMC_25 TSMC_24 VSSI VSSI VDDHD VDDI TSMC_8 
+ S1ALLSVTSW2000X20_nor3_svt_mac_pcell_4 n_totalM=4 n_nfin=6 n_l=16.0n 
+ p_totalM=4 p_nfin=6 p_l=16.0n 
XTSEL_RT TSMC_2 TSMC_33 TSMC_31 TSMC_20 TSMC_21 VDDHD VDDI VSSI TSMC_36 
+ TSMC_37 S1ALLSVTSW2000X20_RESETD_TSEL_M8 
MM22 TSMC_32 TSMC_10 VSSI VSSI nch_svt_mac l=16.0n nfin=5 m=1 
MM21 TSMC_30 TSMC_33 TSMC_24 VSSI nch_svt_mac l=16.0n nfin=4 m=2 
MM16_MIXV_DFTUUU TSMC_34 TSMC_26 VSSI VSSI nch_ulvt_mac l=16.0n nfin=5 
+ m=1 
MM17_MIXV_DFTUUU TSMC_34 TSMC_27 VSSI VSSI nch_ulvt_mac l=16.0n nfin=5 
+ m=1 
MM4 TSMC_1 TSMC_29 VSSI VSSI nch_svt_mac l=20n nfin=6 m=3 
MM1 TSMC_12 TSMC_31 TSMC_24 VSSI nch_svt_mac l=16.0n nfin=4 m=2 
MN7 TSMC_14 TSMC_32 VSSI VSSI nch_svt_mac l=16.0n nfin=7 m=11 
XI686 VSSI VSSI TSMC_38 TSMC_39 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI668_MIXV_DFTUUU VSSI VSSI TSMC_40 TSMC_26 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=3 n_nfin=6 n_l=16.0n 
+ p_totalM=3 p_nfin=6 p_l=16.0n 
XI649 VSSI VSSI TSMC_13 TSMC_41 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI532 VSSI VSSI TSMC_42 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=4 n_nfin=5 n_l=20n p_totalM=4 
+ p_nfin=11 p_l=20n 
XINV0 VSSI VSSI TSMC_3 TSMC_35 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=4 n_l=16.0n 
+ p_totalM=2 p_nfin=4 p_l=16.0n 
XI638 VSSI VSSI TSMC_31 TSMC_33 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI675 VSSI VSSI TSMC_9 TSMC_43 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV5 VSSI VSSI TSMC_3 TSMC_44 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XINV7 VSSI VSSI TSMC_4 TSMC_45 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI634 VSSI VSSI TSMC_46 TSMC_42 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=8 n_l=20n p_totalM=2 
+ p_nfin=8 p_l=20n 
XINV8 VSSI VSSI TSMC_45 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=3 n_l=20n p_totalM=2 
+ p_nfin=4 p_l=20n 
XI642 VSSI VSSI TSMC_6 TSMC_47 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV6 VSSI VSSI TSMC_44 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=5 n_nfin=4 n_l=20n p_totalM=5 
+ p_nfin=6 p_l=20n 
XI654 VSSI VSSI TSMC_48 TSMC_49 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI685 VSSI VSSI TSMC_34 TSMC_38 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XNAND3_MIXV_ULVT TSMC_36 TSMC_37 TSMC_3 VSSI VSSI VDDHD VDDI TSMC_29 
+ S1ALLSVTSW2000X20_nand3_ulvt_mac_pcell_2 n_totalM=2 n_nfin=7 
+ n_l=16.0n p_totalM=2 p_nfin=3 p_l=16.0n 
XI645 TSMC_50 TSMC_15 TSMC_14 VSSI VSSI VDDHD VDDI TSMC_46 
+ S1ALLSVTSW2000X20_nand3_svt_mac_pcell_2 n_totalM=2 n_nfin=5 n_l=20n 
+ p_totalM=2 p_nfin=6 p_l=20n 
XI672_MIXV_DFTUUU TSMC_3 TSMC_41 VSSI VSSI VDDHD VDDI TSMC_40 
+ S1ALLSVTSW2000X20_nand2_ulvt_mac_pcell_0 n_totalM=1 n_nfin=6 n_l=16.0n 
+ p_totalM=1 p_nfin=2 p_l=16.0n 
XI644 TSMC_47 TSMC_1 VSSI VSSI VDDHD VDDI TSMC_30 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
XI674 TSMC_11 TSMC_43 VSSI VSSI VDDI VDDI TSMC_31 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
XI631 TSMC_39 TSMC_24 VSSI VSSI VDDHD VDDI TSMC_32 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=2 n_nfin=5 n_l=16.0n 
+ p_totalM=4 p_nfin=7 p_l=16.0n 
XI615 TSMC_51 TSMC_51 TSMC_51 VSSI VSSI VDDHD VDDI TSMC_52 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI625 TSMC_50 TSMC_50 TSMC_50 VSSI VSSI VDDHD VDDI TSMC_48 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI618 TSMC_52 TSMC_52 TSMC_52 VSSI VSSI VDDHD VDDI TSMC_53 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI621 TSMC_14 TSMC_14 TSMC_14 VSSI VSSI VDDHD VDDI TSMC_51 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI624 TSMC_53 TSMC_53 TSMC_53 VSSI VSSI VDDHD VDDI TSMC_50 
+ S1ALLSVTSW2000X20_tri_svt_mac_pcell_5 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    AWTD_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_AWTD_M8 TSMC_1 TSMC_2 VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:O VDDHD:B VDDI:B VSSI:B 
XI18 VSSI VSSI TSMC_3 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=3 n_nfin=12 n_l=20n p_totalM=5 
+ p_nfin=11 p_l=20n 
XINV1 VSSI VSSI TSMC_1 TSMC_3 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=9 n_l=20n p_totalM=2 
+ p_nfin=7 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    COTH_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_COTH_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 VDDHD 
+ VDDI TSMC_26 TSMC_27 VSSI TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 
*.PININFO  TSMC_1:I TSMC_4:I TSMC_8:I TSMC_9:I TSMC_10:I TSMC_12:I TSMC_13:I 
*.PININFO  TSMC_15:I 
*.PININFO  TSMC_16:I TSMC_17:I TSMC_19:I TSMC_20:I TSMC_22:I TSMC_24:I 
*.PININFO  TSMC_28:I TSMC_33:I 
*.PININFO  TSMC_34:I TSMC_2:O TSMC_3:O TSMC_5:O TSMC_6:O TSMC_7:O TSMC_11:O 
*.PININFO  TSMC_14:O TSMC_18:O TSMC_21:O TSMC_26:O TSMC_27:O TSMC_29:O 
*.PININFO  TSMC_30:O 
*.PININFO  TSMC_32:O TSMC_23:B TSMC_25:B VDDHD:B VDDI:B VSSI:B TSMC_31:B 
XVHILO VDDI TSMC_26 TSMC_27 VSSI S1ALLSVTSW2000X20_VHILO 
XPMCTRL TSMC_10 TSMC_11 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 VDDI VSSI 
+ S1ALLSVTSW2000X20_PMCTRL_M8 
XCKG TSMC_5 TSMC_9 TSMC_12 TSMC_14 TSMC_35 TSMC_22 TSMC_24 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_CKG 
XRESETD TSMC_3 TSMC_5 TSMC_5 TSMC_6 TSMC_7 TSMC_9 TSMC_30 TSMC_35 
+ TSMC_21 TSMC_22 TSMC_24 TSMC_25 VDDHD VDDI VSSI TSMC_28 TSMC_29 TSMC_31 
+ TSMC_32 TSMC_27 TSMC_27 TSMC_13 TSMC_15 TSMC_16 TSMC_33 TSMC_34 
+ S1ALLSVTSW2000X20_RESETD_M8 
XAWTD TSMC_1 TSMC_2 VDDHD VDDI VSSI S1ALLSVTSW2000X20_AWTD_M8 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    ENBUFB_WOBIST
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_ENBUFB_WOBIST TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 VDDHD 
+ VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_13:I TSMC_14:I TSMC_4:O TSMC_5:O 
*.PININFO  TSMC_6:O 
*.PININFO  TSMC_7:O TSMC_8:O TSMC_9:O TSMC_10:O TSMC_11:O TSMC_12:O 
*.PININFO  VDDHD:B VDDI:B VSSI:B 
MM2_MIXV_LS_UUU TSMC_15 TSMC_4 VDDI VDDI pch_ulvt_mac l=20n nfin=2 m=1 
MM1_MIXV_LS_UUU TSMC_16 TSMC_2 TSMC_15 VDDI pch_ulvt_mac l=20n nfin=2 
+ m=1 
MM8 TSMC_10 TSMC_11 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
MM19_MIXV_LS_UUU TSMC_17 TSMC_3 VDDI VDDI pch_ulvt_mac l=16.0n nfin=5 
+ m=2 
MM11 TSMC_18 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=4 m=2 
MM6<1> TSMC_8 TSMC_11 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
MM6<0> TSMC_9 TSMC_11 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
MM7 TSMC_16 TSMC_14 VDDI VDDI pch_svt_mac l=20n nfin=5 m=1 
MM0<1> TSMC_6 TSMC_11 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
MM0<0> TSMC_7 TSMC_11 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=2 
MM10_MIXV_LLS TSMC_11 TSMC_18 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=9 
MM16_MIXV_LS_UUU TSMC_16 TSMC_1 TSMC_17 VDDI pch_ulvt_mac l=16.0n 
+ nfin=5 m=2 
XINV4 VSSI VSSI TSMC_19 TSMC_20 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI148 VSSI VSSI TSMC_4 TSMC_21 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI141 VSSI VSSI TSMC_16 TSMC_4 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=5 n_nfin=4 n_l=20n p_totalM=5 
+ p_nfin=5 p_l=20n 
XI161 VSSI VSSI TSMC_4 TSMC_22 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV7 VSSI VSSI TSMC_23 TSMC_24 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI157 VSSI VSSI TSMC_22 TSMC_12 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI147 VSSI VSSI TSMC_21 TSMC_23 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XINV8 VSSI VSSI TSMC_24 TSMC_25 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
MPD_X1<1> TSMC_8 TSMC_11 VSSI VSSI nch_svt_mac l=20n nfin=12 m=2 
MPD_X1<0> TSMC_9 TSMC_11 VSSI VSSI nch_svt_mac l=20n nfin=12 m=2 
MPD_X2 TSMC_10 TSMC_11 VSSI VSSI nch_svt_mac l=20n nfin=12 m=2 
MM5_MIXV_LS_UUU TSMC_26 TSMC_14 VSSI VSSI nch_ulvt_mac l=20n nfin=2 m=1 
MM17_MIXV_LS_UUU TSMC_16 TSMC_1 TSMC_27 VSSI nch_ulvt_mac l=16.0n 
+ nfin=6 m=2 
MM19_MIXV_LLS TSMC_18 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=3 m=2 
MM18_MIXV_LS_UUU TSMC_27 TSMC_2 TSMC_28 VSSI nch_ulvt_mac l=16.0n 
+ nfin=6 m=2 
MM3_MIXV_LS_UUU TSMC_16 TSMC_3 TSMC_29 VSSI nch_ulvt_mac l=20n nfin=2 
+ m=1 
MM4_MIXV_LS_UUU TSMC_29 TSMC_4 TSMC_26 VSSI nch_ulvt_mac l=20n nfin=2 
+ m=1 
MM21 TSMC_5 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=10 m=14 
MM9 TSMC_11 TSMC_18 VSSI VSSI nch_svt_mac l=20n nfin=3 m=9 
MPD_X0<1> TSMC_6 TSMC_11 VSSI VSSI nch_svt_mac l=20n nfin=12 m=2 
MPD_X0<0> TSMC_7 TSMC_11 VSSI VSSI nch_svt_mac l=20n nfin=12 m=2 
MM20_MIXV_LS_UUU TSMC_28 TSMC_14 VSSI VSSI nch_ulvt_mac l=16.0n nfin=6 
+ m=2 
XI158 TSMC_25 TSMC_25 VSSI VSSI VDDHD VDDI TSMC_19 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DECB1_AND
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DECB1_AND TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI VSSI 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_4:I TSMC_1:O VDDHD:B VDDI:B VSSI:B 
MTN1 TSMC_5 TSMC_4 TSMC_3 VSSI nch_svt_mac l=20n nfin=7 m=1 
MN0 TSMC_1 TSMC_5 VSSI VSSI nch_svt_mac l=20n nfin=12 m=5 
MM3 TSMC_5 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_1 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=12 m=6 
MP5 TSMC_5 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=4 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    CKBUF_M16
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_CKBUF_M16 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI VSSI 
*.PININFO  TSMC_3:I TSMC_4:I TSMC_1:O TSMC_2:O VDDHD:B VDDI:B VSSI:B 
XINV0 VSSI VSSI TSMC_1 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=3 n_nfin=6 n_l=20n p_totalM=3 
+ p_nfin=9 p_l=20n 
MNOR0_N2 TSMC_1 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=6 m=2 
MNOR0_N1 TSMC_1 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=6 m=2 
MNOR0_P2 TSMC_1 TSMC_3 TSMC_5 VDDI pch_svt_mac l=20n nfin=9 m=2 
MNOR0_P1 TSMC_5 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=9 m=2 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    ABUF_WOBIST
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_ABUF_WOBIST TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD 
+ VDDI VSSI 
*.PININFO  TSMC_3:I TSMC_4:I TSMC_5:I TSMC_1:O TSMC_2:O VDDHD:B VDDI:B VSSI:B 
MM21 TSMC_6 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM20 TSMC_2 TSMC_5 TSMC_6 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM19 TSMC_2 TSMC_3 TSMC_8 VSSI nch_svt_mac l=20n nfin=5 m=1 
MM23 TSMC_8 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=5 m=1 
MM27 TSMC_9 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM26 TSMC_2 TSMC_4 TSMC_9 VDDI pch_svt_mac l=20n nfin=2 m=1 
MM29 TSMC_2 TSMC_3 TSMC_10 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM28 TSMC_10 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
XI25 VSSI VSSI TSMC_2 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI54 VSSI VSSI TSMC_2 TSMC_1 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DECB2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DECB2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD VDDI 
+ VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:O TSMC_5:O VDDHD:B VDDI:B VSSI:B 
MM2 TSMC_6 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_6 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_7 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_7 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM0 TSMC_6 TSMC_1 TSMC_8 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM7 TSMC_7 TSMC_2 TSMC_8 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM8 TSMC_8 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
XINV0 VSSI VSSI TSMC_7 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XINV1 VSSI VSSI TSMC_6 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    ABUF_DECB2_WOBIST
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_ABUF_DECB2_WOBIST TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 VDDHD VDDI VSSI TSMC_9 TSMC_10 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:O TSMC_6:O TSMC_7:O 
*.PININFO  TSMC_8:O 
*.PININFO  TSMC_9:O TSMC_10:O VDDHD:B VDDI:B VSSI:B 
XABUF<1> TSMC_10 TSMC_11 TSMC_4 TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ABUF_WOBIST 
XABUF<0> TSMC_9 TSMC_12 TSMC_3 TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ABUF_WOBIST 
XDECB2<1> TSMC_9 TSMC_12 TSMC_11 TSMC_7 TSMC_8 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB2 
XDECB2<0> TSMC_9 TSMC_12 TSMC_10 TSMC_5 TSMC_6 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB2 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DECB4
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DECB4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:O TSMC_7:O 
*.PININFO  TSMC_8:O 
*.PININFO  TSMC_9:O VDDHD:B VDDI:B VSSI:B 
MM15 TSMC_10 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM16 TSMC_10 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM17 TSMC_11 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM18 TSMC_11 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM22 TSMC_11 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM23 TSMC_10 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM24 TSMC_12 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM25 TSMC_13 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM5 TSMC_12 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM4 TSMC_12 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM2 TSMC_13 TSMC_3 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM1 TSMC_13 TSMC_1 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM19 TSMC_14 TSMC_4 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM20 TSMC_10 TSMC_2 TSMC_14 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM21 TSMC_11 TSMC_1 TSMC_14 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM26 TSMC_15 TSMC_5 VSSI VSSI nch_svt_mac l=20n nfin=6 m=1 
MM8 TSMC_16 TSMC_3 TSMC_15 VSSI nch_svt_mac l=20n nfin=3 m=1 
MM7 TSMC_12 TSMC_2 TSMC_16 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM0 TSMC_13 TSMC_1 TSMC_16 VSSI nch_svt_mac l=20n nfin=2 m=1 
XINV3 VSSI VSSI TSMC_10 TSMC_9 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XINV2 VSSI VSSI TSMC_11 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XINV1 VSSI VSSI TSMC_12 TSMC_7 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XINV0 VSSI VSSI TSMC_13 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    ABUF_DECB4_WOBIST
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_ABUF_DECB4_WOBIST TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 VDDHD VDDI VSSI 
+ TSMC_14 TSMC_15 TSMC_16 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:O TSMC_7:O 
*.PININFO  TSMC_8:O 
*.PININFO  TSMC_9:O TSMC_10:O TSMC_11:O TSMC_12:O TSMC_13:O TSMC_14:O TSMC_15:O 
*.PININFO  TSMC_16:O VDDHD:B VDDI:B VSSI:B 
XDECB4<1> TSMC_14 TSMC_17 TSMC_15 TSMC_18 TSMC_19 TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 VDDHD VDDI VSSI S1ALLSVTSW2000X20_DECB4 
XDECB4<0> TSMC_14 TSMC_17 TSMC_15 TSMC_18 TSMC_16 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ VDDHD VDDI VSSI S1ALLSVTSW2000X20_DECB4 
XABUF<2> TSMC_16 TSMC_19 TSMC_5 TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ABUF_WOBIST 
XABUF<0> TSMC_14 TSMC_17 TSMC_3 TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ABUF_WOBIST 
XABUF<1> TSMC_15 TSMC_18 TSMC_4 TSMC_1 TSMC_2 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ABUF_WOBIST 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DECB1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DECB1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 VDDHD 
+ VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_3:O VDDHD:B VDDI:B 
*.PININFO  VSSI:B 
MTN1_MIXV_WAS TSMC_7 TSMC_1 TSMC_8 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2_MIXV_WAS TSMC_8 TSMC_6 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=12 m=2 
MM0_MIXV_WAS TSMC_7 TSMC_2 TSMC_8 VSSI nch_ulvt_mac l=20n nfin=7 m=1 
MN0 TSMC_3 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=12 m=5 
MM1 TSMC_9 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_7 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0 TSMC_3 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=12 m=6 
MP5 TSMC_7 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM2 TSMC_7 TSMC_1 TSMC_9 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DECB1_CKD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DECB1_CKD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_3:O VDDHD:B VDDI:B 
*.PININFO  VSSI:B 
MTN1_MIXV_WAS TSMC_7 TSMC_1 TSMC_8 VSSI nch_ulvt_mac l=20n nfin=3 m=1 
MTN2_MIXV_WAS TSMC_8 TSMC_6 TSMC_5 VSSI nch_ulvt_mac l=20n nfin=12 m=2 
MM0_MIXV_WAS TSMC_7 TSMC_2 TSMC_8 VSSI nch_ulvt_mac l=20n nfin=7 m=1 
MN0_MIXV_DFTUUU TSMC_3 TSMC_7 VSSI VSSI nch_ulvt_mac l=20n nfin=12 m=5 
MM1 TSMC_9 TSMC_2 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MM3 TSMC_7 TSMC_6 VDDHD VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0_MIXV_DFTUUU TSMC_3 TSMC_7 VDDHD VDDI pch_ulvt_mac l=20n nfin=12 m=6 
MP5 TSMC_7 TSMC_4 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM2 TSMC_7 TSMC_1 TSMC_9 VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    ABUF2_WOBIST
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_ABUF2_WOBIST TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VDDHD 
+ VDDI VSSI 
*.PININFO  TSMC_3:I TSMC_4:I TSMC_5:I TSMC_1:O TSMC_2:O VDDHD:B VDDI:B VSSI:B 
MM23 TSMC_6 TSMC_4 VSSI VSSI nch_svt_mac l=20n nfin=5 m=1 
MM21 TSMC_7 TSMC_8 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM20 TSMC_2 TSMC_5 TSMC_7 VSSI nch_svt_mac l=20n nfin=2 m=1 
MM19 TSMC_2 TSMC_3 TSMC_6 VSSI nch_svt_mac l=20n nfin=5 m=1 
MM29 TSMC_2 TSMC_3 TSMC_9 VDDI pch_svt_mac l=20n nfin=5 m=1 
MM28 TSMC_9 TSMC_5 VDDHD VDDI pch_svt_mac l=20n nfin=5 m=1 
MM27 TSMC_10 TSMC_8 VDDHD VDDI pch_svt_mac l=20n nfin=2 m=1 
MM26 TSMC_2 TSMC_4 TSMC_10 VDDI pch_svt_mac l=20n nfin=2 m=1 
XI54 VSSI VSSI TSMC_2 TSMC_1 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI25 VSSI VSSI TSMC_2 TSMC_8 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DECB1_BS_SEG
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DECB1_BS_SEG TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_3:O VDDHD:B VDDI:B 
*.PININFO  VSSI:B 
MTN1_MIXV_WAS TSMC_7 TSMC_1 TSMC_8 VSSI nch_ulvt_mac l=16.0n nfin=3 m=1 
MTN2_MIXV_WAS TSMC_8 TSMC_6 TSMC_5 VSSI nch_ulvt_mac l=16.0n nfin=12 m=2 
MM0_MIXV_WAS TSMC_7 TSMC_2 TSMC_8 VSSI nch_ulvt_mac l=16.0n nfin=7 m=1 
MN0 TSMC_3 TSMC_7 VSSI VSSI nch_svt_mac l=20n nfin=12 m=5 
MM3 TSMC_7 TSMC_6 VDDHD VDDI pch_svt_mac l=16.0n nfin=3 m=1 
MP5 TSMC_7 TSMC_4 VDDHD VDDI pch_svt_mac l=16.0n nfin=5 m=1 
MM2 TSMC_7 TSMC_1 TSMC_9 VDDI pch_svt_mac l=16.0n nfin=3 m=1 
MP0 TSMC_3 TSMC_7 VDDHD VDDI pch_svt_mac l=20n nfin=12 m=6 
MM1 TSMC_9 TSMC_2 VDDHD VDDI pch_svt_mac l=16.0n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    CDEC_M8M16_WOBIST
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_CDEC_M8M16_WOBIST TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 
+ TSMC_61 TSMC_62 TSMC_63 TSMC_64 VDDHD VDDI VSSI TSMC_65 TSMC_66 TSMC_67 
+ TSMC_68 TSMC_69 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I 
*.PININFO  TSMC_8:I 
*.PININFO  TSMC_9:I TSMC_10:I TSMC_11:I TSMC_12:I TSMC_13:I TSMC_14:I TSMC_15:I 
*.PININFO  TSMC_16:I 
*.PININFO  TSMC_19:I TSMC_20:I TSMC_21:I TSMC_22:I TSMC_23:I TSMC_62:I 
*.PININFO  TSMC_63:I TSMC_64:I 
*.PININFO  TSMC_67:I TSMC_17:O TSMC_18:O TSMC_24:O TSMC_25:O TSMC_26:O 
*.PININFO  TSMC_27:O 
*.PININFO  TSMC_28:O TSMC_29:O TSMC_30:O TSMC_31:O TSMC_32:O 
*.PININFO  TSMC_33:O TSMC_34:O TSMC_35:O TSMC_36:O TSMC_37:O 
*.PININFO  TSMC_38:O TSMC_39:O TSMC_40:O TSMC_41:O TSMC_42:O 
*.PININFO  TSMC_43:O TSMC_44:O TSMC_45:O TSMC_46:O TSMC_47:O 
*.PININFO  TSMC_48:O TSMC_49:O TSMC_50:O TSMC_51:O TSMC_52:O 
*.PININFO  TSMC_53:O TSMC_54:O TSMC_55:O TSMC_56:O TSMC_57:O TSMC_58:O 
*.PININFO  TSMC_59:O TSMC_60:O TSMC_61:O TSMC_65:O TSMC_66:O TSMC_68:O 
*.PININFO  TSMC_69:O VDDHD:B VDDI:B 
*.PININFO  VSSI:B 
XCEBBUF TSMC_16 TSMC_70 TSMC_17 TSMC_60 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 
+ TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_64 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ENBUFB_WOBIST 
XIDEC_X2<0> TSMC_40 TSMC_77 TSMC_76 TSMC_80 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X2<1> TSMC_41 TSMC_77 TSMC_76 TSMC_81 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X2<2> TSMC_42 TSMC_77 TSMC_76 TSMC_82 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X2<3> TSMC_43 TSMC_77 TSMC_76 TSMC_83 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<0> TSMC_24 TSMC_77 TSMC_72 TSMC_84 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<1> TSMC_25 TSMC_77 TSMC_72 TSMC_85 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<2> TSMC_26 TSMC_77 TSMC_72 TSMC_86 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<3> TSMC_27 TSMC_77 TSMC_72 TSMC_87 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<4> TSMC_28 TSMC_77 TSMC_73 TSMC_88 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<5> TSMC_29 TSMC_77 TSMC_73 TSMC_89 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<6> TSMC_30 TSMC_77 TSMC_73 TSMC_90 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X0<7> TSMC_31 TSMC_77 TSMC_73 TSMC_91 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<0> TSMC_32 TSMC_77 TSMC_74 TSMC_92 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<1> TSMC_33 TSMC_77 TSMC_74 TSMC_93 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<2> TSMC_34 TSMC_77 TSMC_74 TSMC_94 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<3> TSMC_35 TSMC_77 TSMC_74 TSMC_95 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<4> TSMC_36 TSMC_77 TSMC_75 TSMC_96 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<5> TSMC_37 TSMC_77 TSMC_75 TSMC_97 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<6> TSMC_38 TSMC_77 TSMC_75 TSMC_98 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XIDEC_X1<7> TSMC_39 TSMC_77 TSMC_75 TSMC_99 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_AND 
XCKBUF TSMC_70 TSMC_17 TSMC_19 TSMC_23 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_CKBUF_M16 
XABUF_PDEC_X2 TSMC_70 TSMC_17 TSMC_7 TSMC_8 TSMC_80 TSMC_81 TSMC_82 TSMC_83 
+ VDDHD VDDI VSSI TSMC_100 TSMC_101 
+ S1ALLSVTSW2000X20_ABUF_DECB2_WOBIST 
XABUF_PDEC_Y TSMC_70 TSMC_17 TSMC_12 TSMC_13 TSMC_14 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 VDDHD VDDI VSSI 
+ TSMC_110 TSMC_111 TSMC_112 S1ALLSVTSW2000X20_ABUF_DECB4_WOBIST 
XABUF_PDEC_X0 TSMC_70 TSMC_17 TSMC_1 TSMC_2 TSMC_3 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 VDDHD VDDI VSSI TSMC_113 
+ TSMC_114 TSMC_115 S1ALLSVTSW2000X20_ABUF_DECB4_WOBIST 
XABUF_PDEC_X1 TSMC_70 TSMC_17 TSMC_4 TSMC_5 TSMC_6 TSMC_92 TSMC_93 TSMC_94 
+ TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 VDDHD VDDI VSSI TSMC_116 
+ TSMC_117 TSMC_118 S1ALLSVTSW2000X20_ABUF_DECB4_WOBIST 
XABUF_PDEC_X3 TSMC_70 TSMC_17 TSMC_9 TSMC_10 TSMC_11 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 VDDHD VDDI VSSI 
+ TSMC_127 TSMC_128 TSMC_129 S1ALLSVTSW2000X20_ABUF_DECB4_WOBIST 
XIDEC_WE TSMC_20 TSMC_23 TSMC_65 TSMC_77 TSMC_71 TSMC_66 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_YL<0> TSMC_20 TSMC_23 TSMC_68 TSMC_77 TSMC_71 TSMC_130 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_YL<1> TSMC_20 TSMC_23 TSMC_69 TSMC_77 TSMC_71 TSMC_131 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_RE TSMC_20 TSMC_23 TSMC_61 TSMC_77 TSMC_71 TSMC_132 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<0> TSMC_20 TSMC_23 TSMC_52 TSMC_77 TSMC_71 TSMC_102 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<1> TSMC_20 TSMC_23 TSMC_53 TSMC_77 TSMC_71 TSMC_103 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<2> TSMC_20 TSMC_23 TSMC_54 TSMC_77 TSMC_71 TSMC_104 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<3> TSMC_20 TSMC_23 TSMC_55 TSMC_77 TSMC_71 TSMC_105 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<4> TSMC_20 TSMC_23 TSMC_56 TSMC_77 TSMC_71 TSMC_106 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<5> TSMC_20 TSMC_23 TSMC_57 TSMC_77 TSMC_71 TSMC_107 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<6> TSMC_20 TSMC_23 TSMC_58 TSMC_77 TSMC_71 TSMC_108 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_Y<7> TSMC_20 TSMC_23 TSMC_59 TSMC_77 TSMC_71 TSMC_109 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1 
XIDEC_CKD TSMC_21 TSMC_23 TSMC_18 TSMC_78 TSMC_71 TSMC_66 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_DECB1_CKD 
XABUF_Y<3> TSMC_130 TSMC_133 TSMC_15 TSMC_70 TSMC_17 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ABUF2_WOBIST 
XWEBBUF TSMC_66 TSMC_134 TSMC_67 TSMC_70 TSMC_17 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_ABUF2_WOBIST 
XI27 VSSI VSSI TSMC_130 TSMC_131 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XI303 VSSI VSSI TSMC_66 TSMC_132 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XIDEC_X3<0> TSMC_19 TSMC_23 TSMC_44 TSMC_60 TSMC_71 TSMC_119 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
XIDEC_X3<1> TSMC_19 TSMC_23 TSMC_45 TSMC_60 TSMC_71 TSMC_120 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
XIDEC_X3<2> TSMC_19 TSMC_23 TSMC_46 TSMC_60 TSMC_71 TSMC_121 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
XIDEC_X3<3> TSMC_19 TSMC_23 TSMC_47 TSMC_60 TSMC_71 TSMC_122 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
XIDEC_X3<4> TSMC_19 TSMC_23 TSMC_48 TSMC_60 TSMC_71 TSMC_123 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
XIDEC_X3<5> TSMC_19 TSMC_23 TSMC_49 TSMC_60 TSMC_71 TSMC_124 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
XIDEC_X3<6> TSMC_19 TSMC_23 TSMC_50 TSMC_60 TSMC_71 TSMC_125 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
XIDEC_X3<7> TSMC_19 TSMC_23 TSMC_51 TSMC_60 TSMC_71 TSMC_126 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_DECB1_BS_SEG 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    CNT_CORE_M8_RWA_WOBIST
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_CNT_CORE_M8_RWA_WOBIST TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 VDDHD 
+ VDDI TSMC_78 TSMC_79 VSSI TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_8:I 
*.PININFO  TSMC_9:I 
*.PININFO  TSMC_10:I TSMC_11:I TSMC_12:I TSMC_13:I TSMC_14:I TSMC_15:I 
*.PININFO  TSMC_16:I TSMC_17:I 
*.PININFO  TSMC_19:I TSMC_21:I TSMC_22:I TSMC_59:I TSMC_62:I TSMC_64:I 
*.PININFO  TSMC_65:I 
*.PININFO  TSMC_66:I TSMC_67:I TSMC_68:I TSMC_70:I TSMC_71:I TSMC_72:I 
*.PININFO  TSMC_75:I TSMC_76:I 
*.PININFO  TSMC_80:I TSMC_81:I TSMC_83:I TSMC_88:I TSMC_89:I TSMC_2:O 
*.PININFO  TSMC_18:O TSMC_20:O TSMC_23:O TSMC_24:O TSMC_25:O TSMC_26:O 
*.PININFO  TSMC_27:O TSMC_28:O TSMC_29:O TSMC_30:O TSMC_31:O 
*.PININFO  TSMC_32:O TSMC_33:O TSMC_34:O TSMC_35:O TSMC_36:O 
*.PININFO  TSMC_37:O TSMC_38:O TSMC_39:O TSMC_40:O TSMC_41:O 
*.PININFO  TSMC_42:O TSMC_43:O TSMC_44:O TSMC_45:O TSMC_46:O 
*.PININFO  TSMC_47:O TSMC_48:O TSMC_49:O TSMC_50:O TSMC_51:O 
*.PININFO  TSMC_52:O TSMC_53:O TSMC_54:O TSMC_55:O TSMC_56:O TSMC_57:O 
*.PININFO  TSMC_58:O TSMC_60:O TSMC_61:O TSMC_63:O TSMC_69:O TSMC_73:O 
*.PININFO  TSMC_78:O TSMC_79:O 
*.PININFO  TSMC_82:O TSMC_84:O TSMC_85:O TSMC_87:O TSMC_90:O TSMC_91:O 
*.PININFO  TSMC_74:B 
*.PININFO  TSMC_77:B VDDHD:B VDDI:B VSSI:B TSMC_86:B 
XMCTRL_RWA TSMC_61 TSMC_72 TSMC_76 VDDHD VDDI VSSI TSMC_80 TSMC_81 
+ TSMC_20 S1ALLSVTSW2000X20_MCTRL_RWA_M8 
XCOTHERS TSMC_1 TSMC_2 TSMC_18 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_21 TSMC_22 
+ TSMC_59 TSMC_60 TSMC_96 TSMC_62 TSMC_97 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_73 TSMC_72 TSMC_74 TSMC_75 TSMC_77 VDDHD 
+ VDDI TSMC_78 TSMC_79 VSSI TSMC_98 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_89 S1ALLSVTSW2000X20_COTH_M8 
XCDEC TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 
+ TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_19 TSMC_92 TSMC_20 
+ TSMC_93 TSMC_94 TSMC_95 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_96 TSMC_63 TSMC_64 TSMC_65 TSMC_97 VDDHD VDDI VSSI 
+ TSMC_82 TSMC_98 TSMC_83 TSMC_90 TSMC_91 
+ S1ALLSVTSW2000X20_CDEC_M8M16_WOBIST 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    TM_BUF_DSLP_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_TM_BUF_DSLP_M8 TSMC_1 TSMC_2 TSMC_3 VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_3:I VDDI:I VSSI:I TSMC_2:O 
XI2 VSSI VSSI TSMC_4 TSMC_2 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI4 VSSI VSSI TSMC_3 TSMC_5 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI3 TSMC_1 TSMC_5 VSSI VSSI VDDI VDDI TSMC_4 
+ S1ALLSVTSW2000X20_nand2_svt_mac_pcell_0 n_totalM=1 n_nfin=2 n_l=20n 
+ p_totalM=1 p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    CNT_M8_IOX4
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_CNT_M8_IOX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 VDDHD VDDI TSMC_117 TSMC_118 VSSI TSMC_119 
+ TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 
+ TSMC_128 TSMC_129 TSMC_130 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_6:I TSMC_7:I TSMC_8:I 
*.PININFO  TSMC_9:I 
*.PININFO  TSMC_10:I TSMC_11:I TSMC_12:I TSMC_13:I TSMC_14:I TSMC_15:I 
*.PININFO  TSMC_16:I TSMC_17:I 
*.PININFO  TSMC_19:I TSMC_20:I TSMC_21:I TSMC_22:I TSMC_23:I TSMC_25:I 
*.PININFO  TSMC_26:I TSMC_63:I 
*.PININFO  TSMC_66:I TSMC_67:I TSMC_69:I TSMC_70:I TSMC_71:I TSMC_72:I 
*.PININFO  TSMC_90:I 
*.PININFO  TSMC_96:I TSMC_97:I TSMC_98:I TSMC_99:I TSMC_100:I TSMC_102:I 
*.PININFO  TSMC_104:I 
*.PININFO  TSMC_107:I TSMC_108:I TSMC_112:I TSMC_113:I TSMC_114:I TSMC_119:I 
*.PININFO  TSMC_120:I TSMC_122:I TSMC_127:I TSMC_128:I TSMC_64:O TSMC_65:O 
*.PININFO  TSMC_81:O TSMC_82:O TSMC_83:O TSMC_84:O TSMC_85:O TSMC_86:O 
*.PININFO  TSMC_87:O TSMC_88:O 
*.PININFO  TSMC_91:O TSMC_92:O TSMC_93:O TSMC_94:O TSMC_105:O TSMC_106:O 
*.PININFO  TSMC_115:O TSMC_2:B 
*.PININFO  TSMC_18:B TSMC_24:B TSMC_27:B TSMC_28:B TSMC_29:B TSMC_30:B 
*.PININFO  TSMC_31:B TSMC_32:B TSMC_33:B TSMC_34:B TSMC_35:B 
*.PININFO  TSMC_36:B TSMC_37:B TSMC_38:B TSMC_39:B TSMC_40:B 
*.PININFO  TSMC_41:B TSMC_42:B TSMC_43:B TSMC_44:B TSMC_45:B 
*.PININFO  TSMC_46:B TSMC_47:B TSMC_48:B TSMC_49:B TSMC_50:B 
*.PININFO  TSMC_51:B TSMC_52:B TSMC_53:B TSMC_54:B TSMC_55:B 
*.PININFO  TSMC_56:B TSMC_57:B TSMC_58:B TSMC_59:B TSMC_60:B TSMC_61:B 
*.PININFO  TSMC_62:B TSMC_68:B TSMC_73:B TSMC_74:B TSMC_75:B TSMC_76:B 
*.PININFO  TSMC_77:B 
*.PININFO  TSMC_78:B TSMC_79:B TSMC_80:B TSMC_89:B TSMC_95:B TSMC_101:B 
*.PININFO  TSMC_103:B 
*.PININFO  TSMC_109:B TSMC_110:B TSMC_111:B TSMC_116:B VDDHD:B VDDI:B 
*.PININFO  TSMC_117:B TSMC_118:B 
*.PININFO  VSSI:B TSMC_121:B TSMC_123:B TSMC_124:B TSMC_125:B TSMC_126:B 
*.PININFO  TSMC_129:B TSMC_130:B 
MM4<0> TSMC_35 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4<1> TSMC_36 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4<2> TSMC_37 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4<3> TSMC_38 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4<4> TSMC_39 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4<5> TSMC_40 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4<6> TSMC_41 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM4<7> TSMC_42 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<0> TSMC_27 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<1> TSMC_28 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<2> TSMC_29 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<3> TSMC_30 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<4> TSMC_31 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<5> TSMC_32 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<6> TSMC_33 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MX0_PD<7> TSMC_34 TSMC_106 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
XIO_L TSMC_2 TSMC_21 TSMC_24 TSMC_71 TSMC_79 TSMC_77 TSMC_87 TSMC_85 TSMC_93 
+ TSMC_106 VDDHD VDDI VSSI TSMC_124 TSMC_126 
+ S1ALLSVTSW2000X20_IO_INV_NM 
XIO_R TSMC_2 TSMC_22 TSMC_24 TSMC_72 TSMC_80 TSMC_78 TSMC_88 TSMC_86 TSMC_94 
+ TSMC_106 VDDHD VDDI VSSI TSMC_124 TSMC_126 
+ S1ALLSVTSW2000X20_IO_INV_NM 
XIO_RR TSMC_2 TSMC_20 TSMC_24 TSMC_70 TSMC_74 TSMC_76 TSMC_82 TSMC_84 TSMC_92 
+ TSMC_106 VDDHD VDDI VSSI TSMC_124 TSMC_126 
+ S1ALLSVTSW2000X20_IO_INV_NM 
XIO_LL TSMC_2 TSMC_19 TSMC_24 TSMC_69 TSMC_73 TSMC_75 TSMC_81 TSMC_83 TSMC_91 
+ TSMC_106 VDDHD VDDI VSSI TSMC_124 TSMC_126 
+ S1ALLSVTSW2000X20_IO_INV_NM 
XI72_MIXV_UHD TSMC_103 TSMC_103 VSSI VSSI VDDI VDDI TSMC_131 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
MVDDHD_GG_MIXV_HD4 VDDHD TSMC_105 VDDI VDDI pch_svt_mac l=20n nfin=10 
+ m=140 
MVDDHD_GG_MIXV_HD VDDHD TSMC_103 VDDI VDDI pch_svt_mac l=20n nfin=10 
+ m=40 
MVDDHD_GG_MIXV_HD2 VDDHD TSMC_103 VDDI VDDI pch_svt_mac l=20n nfin=12 
+ m=10 
MVDDHD_GG_MIXV_HD3 VDDHD TSMC_103 VDDI VDDI pch_svt_mac l=20n nfin=8 
+ m=7 
XTMWAS_CAP_BUF TSMC_114 TSMC_115 TSMC_106 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_TM_BUF 
XCNT TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 
+ TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 
+ TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 
+ TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_68 TSMC_89 TSMC_90 TSMC_95 TSMC_96 TSMC_97 TSMC_98 
+ TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_108 TSMC_106 TSMC_103 
+ TSMC_111 TSMC_112 TSMC_113 TSMC_116 VDDHD VDDI TSMC_117 TSMC_118 VSSI 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ S1ALLSVTSW2000X20_CNT_CORE_M8_RWA_WOBIST 
XI10 VSSI VSSI TSMC_131 TSMC_105 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=3 n_nfin=11 n_l=20n p_totalM=1 
+ p_nfin=11 p_l=20n 
XI11 VSSI VSSI TSMC_131 TSMC_106 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=5 n_nfin=7 n_l=20n p_totalM=1 
+ p_nfin=11 p_l=20n 
XDSLPSEL_BUF<0> TSMC_66 TSMC_64 TSMC_100 VDDI VSSI 
+ S1ALLSVTSW2000X20_TM_BUF_DSLP_M8 
XDSLPSEL_BUF<1> TSMC_67 TSMC_65 TSMC_100 VDDI VSSI 
+ S1ALLSVTSW2000X20_TM_BUF_DSLP_M8 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    DIO
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_DIO TSMC_1 TSMC_2 
*.PININFO  TSMC_1:B TSMC_2:B 
XD7 TSMC_2 TSMC_1 ndio_mac nfin=2 l=200n m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    BUF_IO2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_BUF_IO2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:O TSMC_4:O VDDHD:B VDDI:B VSSI:B 
XI364<1> VSSI VSSI TSMC_5 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI364<0> VSSI VSSI TSMC_2 TSMC_5 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI0<1> VSSI VSSI TSMC_6 TSMC_3 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI0<0> VSSI VSSI TSMC_1 TSMC_6 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    VLO
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_VLO VDDI TSMC_1 TSMC_2 VSSI 
*.PININFO  TSMC_1:O TSMC_2:O VDDI:B VSSI:B 
MN3 VSSI TSMC_3 TSMC_4 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN0 VSSI TSMC_4 TSMC_4 VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1 VSSI TSMC_3 TSMC_2 VSSI nch_svt_mac l=20n nfin=6 m=2 
MP7 TSMC_3 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP2 TSMC_1 TSMC_4 VDDI VDDI pch_svt_mac l=20n nfin=12 m=1 
MP0 TSMC_3 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    IO_M8B
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_IO_M8B TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 VDDHD VDDI VSSI TSMC_12 TSMC_13 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_11:I TSMC_12:I TSMC_13:I 
*.PININFO  TSMC_7:O TSMC_8:O 
*.PININFO  TSMC_10:O TSMC_5:B TSMC_6:B TSMC_9:B VDDHD:B VDDI:B VSSI:B 
MP1_MIXV_HD VDDHD TSMC_9 VDDI VDDI pch_svt_mac l=20n nfin=10 m=11 
XIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_10 TSMC_11 
+ VDDHD VDDI VSSI TSMC_12 TSMC_13 S1ALLSVTSW2000X20_IO_INV_NM 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    LCTRL_PM_S
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_LCTRL_PM_S TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_4:I TSMC_5:I TSMC_2:O TSMC_3:O TSMC_6:O VDDI:B VSSI:B 
XI255 TSMC_5 TSMC_1 TSMC_4 VSSI VSSI VDDI VDDI TSMC_7 
+ S1ALLSVTSW2000X20_nor3_svt_mac_pcell_4 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI257 VSSI VSSI TSMC_5 TSMC_8 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI232 VSSI VSSI TSMC_8 TSMC_2 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=7 n_l=20n p_totalM=1 
+ p_nfin=7 p_l=20n 
XI256 VSSI VSSI TSMC_7 TSMC_6 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    LCTRL_BUF_S
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_LCTRL_BUF_S TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VDDAI VDDI TSMC_7 TSMC_8 VSSI 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_7:O TSMC_8:O TSMC_3:B TSMC_4:B 
*.PININFO  TSMC_5:B TSMC_6:B VDDAI:B VDDI:B VSSI:B 
MM59 TSMC_5 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=5 m=1 
MM1 TSMC_4 TSMC_6 VDDI VDDI pch_svt_mac l=20n nfin=10 m=2 
MM56 TSMC_6 TSMC_5 VDDI VDDI pch_svt_mac l=20n nfin=10 m=1 
MM0 TSMC_4 TSMC_6 VSSI VSSI nch_svt_mac l=20n nfin=10 m=2 
MM46 TSMC_5 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=5 m=1 
MM52 TSMC_6 TSMC_5 VSSI VSSI nch_svt_mac l=20n nfin=10 m=1 
XVHILO VDDI TSMC_7 TSMC_8 VSSI S1ALLSVTSW2000X20_VLO 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    TRKBL_ISO_X2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_TRKBL_ISO_X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
*.PININFO  TSMC_9:B 
Mpg11 TSMC_1 TSMC_2 TSMC_10 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd11 TSMC_10 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_11 TSMC_10 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg21 TSMC_12 TSMC_7 TSMC_11 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_13 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_14 TSMC_13 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_13 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_12 TSMC_8 TSMC_14 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
MM0 TSMC_15 TSMC_10 TSMC_9 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu11 TSMC_10 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_13 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    TRKBL_OFF_X2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_TRKBL_OFF_X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
Mpg11 TSMC_1 TSMC_4 TSMC_9 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd11 TSMC_9 TSMC_10 TSMC_11 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_4 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg21 TSMC_12 TSMC_5 TSMC_10 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_13 TSMC_14 TSMC_11 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_14 TSMC_13 TSMC_4 TSMC_4 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_4 TSMC_13 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_12 TSMC_6 TSMC_14 TSMC_4 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpu11 TSMC_9 TSMC_10 TSMC_3 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_13 TSMC_14 TSMC_3 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu21 TSMC_10 TSMC_9 TSMC_8 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu20 TSMC_14 TSMC_13 TSMC_7 TSMC_2 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    MCB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_MCB TSMC_1 TSMC_2 VDDAI VDDI VSSI TSMC_3 
*.PININFO  TSMC_1:B TSMC_2:B VDDAI:B VDDI:B VSSI:B TSMC_3:B 
MM4 TSMC_4 TSMC_5 VDDAI VDDI pchpu_hcsr_mac l=20n nfin=1 m=1 
MM6 TSMC_5 TSMC_4 VDDAI VDDI pchpu_hcsr_mac l=20n nfin=1 m=1 
MM0 TSMC_1 TSMC_3 TSMC_5 VSSI nchpg_hcsr_mac l=20n nfin=2 m=1 
MM5 TSMC_2 TSMC_3 TSMC_4 VSSI nchpg_hcsr_mac l=20n nfin=2 m=1 
MM1 TSMC_5 TSMC_4 VSSI VSSI nchpd_hcsr_mac l=20n nfin=2 m=1 
MM2 TSMC_4 TSMC_5 VSSI VSSI nchpd_hcsr_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    TRKBL_ON_X2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_TRKBL_ON_X2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
Mpg11 TSMC_1 TSMC_2 TSMC_9 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd11 TSMC_9 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd21 TSMC_10 TSMC_9 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg21 TSMC_11 TSMC_7 TSMC_10 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpd10 TSMC_12 TSMC_5 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpd20 TSMC_13 TSMC_12 TSMC_6 TSMC_6 nchpd_hcsr_mac l=20n nfin=2 m=1 
Mpg10 TSMC_1 TSMC_3 TSMC_12 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpg20 TSMC_11 TSMC_8 TSMC_13 TSMC_6 nchpg_hcsr_mac l=20n nfin=2 m=1 
Mpu11 TSMC_9 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
Mpu10 TSMC_12 TSMC_5 TSMC_5 TSMC_4 pchpu_hcsr_mac l=20n nfin=1 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    MCB_2X8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_MCB_2X8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_21 TSMC_22 
*.PININFO  TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B TSMC_7:B 
*.PININFO  TSMC_8:B 
*.PININFO  TSMC_9:B TSMC_10:B TSMC_11:B TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B 
*.PININFO  TSMC_16:B TSMC_17:B TSMC_18:B TSMC_19:B TSMC_20:B VDDAI:B VDDI:B 
*.PININFO  VSSI:B TSMC_21:B 
*.PININFO  TSMC_22:B 
XMCB_1<0> TSMC_1 TSMC_9 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_1<1> TSMC_2 TSMC_10 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_1<2> TSMC_3 TSMC_11 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_1<3> TSMC_4 TSMC_12 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_1<4> TSMC_5 TSMC_13 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_1<5> TSMC_6 TSMC_14 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_1<6> TSMC_7 TSMC_15 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_1<7> TSMC_8 TSMC_16 VDDAI VDDI VSSI TSMC_22 S1ALLSVTSW2000X20_MCB 
XMCB_0<0> TSMC_1 TSMC_9 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
XMCB_0<1> TSMC_2 TSMC_10 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
XMCB_0<2> TSMC_3 TSMC_11 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
XMCB_0<3> TSMC_4 TSMC_12 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
XMCB_0<4> TSMC_5 TSMC_13 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
XMCB_0<5> TSMC_6 TSMC_14 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
XMCB_0<6> TSMC_7 TSMC_15 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
XMCB_0<7> TSMC_8 TSMC_16 VDDAI VDDI VSSI TSMC_21 S1ALLSVTSW2000X20_MCB 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    TOP_EDGE2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_TOP_EDGE2 VDDHD VDDI VSSI TSMC_1 TSMC_2 
*.PININFO  VDDHD:B VDDI:B VSSI:B TSMC_1:B TSMC_2:B 
XI56 VSSI VSSI TSMC_3 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=8 n_l=20n p_totalM=2 
+ p_nfin=10 p_l=20n 
XI59 VSSI VSSI TSMC_3 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=8 n_l=20n p_totalM=2 
+ p_nfin=10 p_l=20n 
XI58 VSSI VSSI TSMC_3 TSMC_4 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=8 n_l=20n p_totalM=2 
+ p_nfin=10 p_l=20n 
XI57 VSSI VSSI TSMC_3 TSMC_2 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=8 n_l=20n p_totalM=2 
+ p_nfin=10 p_l=20n 
XI55 VSSI VSSI TSMC_1 TSMC_3 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=7 n_l=20n p_totalM=1 
+ p_nfin=10 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WOBIST_IO2
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WOBIST_IO2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ VSSI 
*.PININFO  TSMC_2:I TSMC_3:I TSMC_1:O TSMC_4:O TSMC_5:B TSMC_6:B VSSI:B 
MM32 TSMC_1 TSMC_2 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM29 TSMC_4 TSMC_3 VSSI VSSI nch_svt_mac l=20n nfin=2 m=1 
MM35 TSMC_1 TSMC_2 TSMC_6 TSMC_5 pch_svt_mac l=20n nfin=2 m=1 
MM25 TSMC_4 TSMC_3 TSMC_6 TSMC_5 pch_svt_mac l=20n nfin=2 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WOBIST_WOLS_IO
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WOBIST_WOLS_IO TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI 
+ VSSI 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_2:O TSMC_4:O VDDHD:B VDDI:B VSSI:B 
XBIST_IO TSMC_5 TSMC_1 TSMC_3 TSMC_6 VDDI VDDHD VSSI 
+ S1ALLSVTSW2000X20_WOBIST_IO2 
XBUF_IO TSMC_5 TSMC_6 TSMC_2 TSMC_4 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_BUF_IO2 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WOBIST_WOLS_IO_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_3:I TSMC_5:I TSMC_2:O TSMC_4:O TSMC_6:B VDDHD:B VDDI:B 
*.PININFO  VSSI:B 
XIO_INTERFACE TSMC_1 TSMC_2 TSMC_3 TSMC_4 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WOBIST_ABUF
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WOBIST_ABUF TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 VSSI 
*.PININFO  TSMC_1:I TSMC_2:O TSMC_3:O TSMC_4:B TSMC_5:B VSSI:B 
MM16 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=4 m=1 
MM30 TSMC_2 TSMC_1 TSMC_4 TSMC_5 pch_svt_mac l=20n nfin=4 m=1 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WOBIST_WOLS_ABUF
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF TSMC_1 TSMC_2 VDDHD VDDI VSSI 
*.PININFO  TSMC_1:I TSMC_2:O VDDHD:B VDDI:B VSSI:B 
XBIST_IO TSMC_1 TSMC_2 TSMC_3 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_ABUF 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WOBIST_WOLS_CNT_M8_IOX4
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WOBIST_WOLS_CNT_M8_IOX4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 VDDHD 
+ VDDI TSMC_33 TSMC_34 VSSI TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 
+ TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 
+ TSMC_68 TSMC_69 TSMC_70 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_8:I TSMC_9:I TSMC_10:I TSMC_12:I 
*.PININFO  TSMC_14:I 
*.PININFO  TSMC_15:I TSMC_16:I TSMC_21:I TSMC_22:I TSMC_27:I TSMC_28:I 
*.PININFO  TSMC_29:I TSMC_30:I TSMC_31:I 
*.PININFO  TSMC_32:I TSMC_35:I TSMC_36:I TSMC_37:I TSMC_39:I TSMC_40:I 
*.PININFO  TSMC_52:I 
*.PININFO  TSMC_53:I TSMC_54:I TSMC_55:I TSMC_56:I TSMC_57:I TSMC_58:I 
*.PININFO  TSMC_59:I TSMC_60:I TSMC_61:I 
*.PININFO  TSMC_62:I TSMC_67:I TSMC_68:I TSMC_69:I TSMC_70:I TSMC_4:O TSMC_5:O 
*.PININFO  TSMC_6:O 
*.PININFO  TSMC_7:O TSMC_11:O TSMC_13:O TSMC_17:O TSMC_18:O TSMC_19:O TSMC_20:O 
*.PININFO  TSMC_33:O 
*.PININFO  TSMC_34:O TSMC_38:O TSMC_41:O TSMC_42:O TSMC_43:O TSMC_44:O 
*.PININFO  TSMC_45:O 
*.PININFO  TSMC_46:O TSMC_47:O TSMC_48:O TSMC_49:O TSMC_50:O TSMC_51:O 
*.PININFO  TSMC_63:O 
*.PININFO  TSMC_64:O TSMC_65:O TSMC_66:O TSMC_23:B TSMC_24:B TSMC_25:B 
*.PININFO  TSMC_26:B VDDHD:B 
*.PININFO  VDDI:B VSSI:B 
XVHILO_VDD_OUT VDDI TSMC_33 TSMC_34 VSSI S1ALLSVTSW2000X20_VHILO 
XBIST_LS_CEB TSMC_10 TSMC_11 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_WEB TSMC_37 TSMC_38 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AY<0> TSMC_67 TSMC_63 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AY<1> TSMC_68 TSMC_64 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AY<2> TSMC_69 TSMC_65 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AY<3> TSMC_70 TSMC_66 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<0> TSMC_52 TSMC_41 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<1> TSMC_53 TSMC_42 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<2> TSMC_54 TSMC_43 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<3> TSMC_55 TSMC_44 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<4> TSMC_56 TSMC_45 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<5> TSMC_57 TSMC_46 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<6> TSMC_58 TSMC_47 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<7> TSMC_59 TSMC_48 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<8> TSMC_60 TSMC_49 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<9> TSMC_61 TSMC_50 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XBIST_LS_ABUF_AX<10> TSMC_62 TSMC_51 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_ABUF 
XINV1 VSSI VSSI TSMC_71 TSMC_13 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=4 n_nfin=5 n_l=16.0n 
+ p_totalM=4 p_nfin=5 p_l=16.0n 
XINV0 VSSI VSSI TSMC_12 TSMC_71 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=5 n_l=16.0n 
+ p_totalM=2 p_nfin=5 p_l=16.0n 
XBIST_LS_IO<1> TSMC_3 TSMC_5 TSMC_15 TSMC_18 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO 
XBIST_LS_IO_R TSMC_9 TSMC_7 TSMC_22 TSMC_20 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO 
XBIST_LS_IO_L TSMC_8 TSMC_6 TSMC_21 TSMC_19 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO 
XBIST_LS_IO<0> TSMC_2 TSMC_4 TSMC_14 TSMC_17 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    IO_M8
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_IO_M8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 VDDHD VDDI VSSI 
+ TSMC_15 TSMC_16 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_9:I TSMC_10:I TSMC_13:I 
*.PININFO  TSMC_15:I 
*.PININFO  TSMC_16:I TSMC_7:O TSMC_8:O TSMC_11:O TSMC_12:O TSMC_14:O TSMC_5:B 
*.PININFO  TSMC_6:B VDDHD:B 
*.PININFO  VDDI:B VSSI:B 
XI159 VSSI VSSI TSMC_17 TSMC_11 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=12 n_nfin=10 n_l=20n 
+ p_totalM=12 p_nfin=10 p_l=20n 
XI161 VSSI VSSI TSMC_13 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI160 VSSI VSSI TSMC_18 TSMC_14 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=3 n_nfin=6 n_l=20n p_totalM=2 
+ p_nfin=6 p_l=20n 
XIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_12 TSMC_14 
+ VDDHD VDDI VSSI TSMC_15 TSMC_16 S1ALLSVTSW2000X20_IO_INV_NM 
MP1_MIXV_HD VDDHD TSMC_11 VDDI VDDI pch_svt_mac l=20n nfin=10 m=11 
XI1 TSMC_9 TSMC_10 VSSI VSSI VDDI VDDI TSMC_17 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=9 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    YPASS_M8_NOSD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_YPASS_M8_NOSD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 VDDAI VDDI VSSI TSMC_22 
+ TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 
+ TSMC_32 
*.PININFO  TSMC_17:I TSMC_21:I TSMC_23:I TSMC_25:I TSMC_26:I TSMC_27:I 
*.PININFO  TSMC_28:I TSMC_29:I TSMC_30:I 
*.PININFO  TSMC_31:I TSMC_32:I TSMC_18:O TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B 
*.PININFO  TSMC_5:B 
*.PININFO  TSMC_6:B TSMC_7:B TSMC_8:B TSMC_9:B TSMC_10:B TSMC_11:B TSMC_12:B 
*.PININFO  TSMC_13:B 
*.PININFO  TSMC_14:B TSMC_15:B TSMC_16:B TSMC_19:B TSMC_20:B VDDAI:B VDDI:B 
*.PININFO  VSSI:B TSMC_22:B TSMC_24:B 
MINV0_M1_MIXV_DFTUUU TSMC_18 TSMC_17 VDDI VDDI pch_ulvt_mac l=20n 
+ nfin=3 m=1 
MM0_MIXV_USD TSMC_19 TSMC_18 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP17<0> TSMC_33 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP17<1> TSMC_34 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP17<2> TSMC_35 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP17<3> TSMC_36 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP17<4> TSMC_37 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP17<5> TSMC_38 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP17<6> TSMC_39 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP17<7> TSMC_40 TSMC_21 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP10_MIXV_USD<0> TSMC_20 TSMC_33 TSMC_9 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP10_MIXV_USD<1> TSMC_20 TSMC_34 TSMC_10 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP10_MIXV_USD<2> TSMC_20 TSMC_35 TSMC_11 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP10_MIXV_USD<3> TSMC_20 TSMC_36 TSMC_12 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP10_MIXV_USD<4> TSMC_20 TSMC_37 TSMC_13 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP10_MIXV_USD<5> TSMC_20 TSMC_38 TSMC_14 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP10_MIXV_USD<6> TSMC_20 TSMC_39 TSMC_15 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP10_MIXV_USD<7> TSMC_20 TSMC_40 TSMC_16 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP3_MIXV_USD TSMC_20 TSMC_18 VDDI VDDI pch_svt_mac l=20n nfin=3 m=1 
MP0_MIXV_USD<0> TSMC_19 TSMC_33 TSMC_1 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP0_MIXV_USD<1> TSMC_19 TSMC_34 TSMC_2 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP0_MIXV_USD<2> TSMC_19 TSMC_35 TSMC_3 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP0_MIXV_USD<3> TSMC_19 TSMC_36 TSMC_4 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP0_MIXV_USD<4> TSMC_19 TSMC_37 TSMC_5 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP0_MIXV_USD<5> TSMC_19 TSMC_38 TSMC_6 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP0_MIXV_USD<6> TSMC_19 TSMC_39 TSMC_7 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP0_MIXV_USD<7> TSMC_19 TSMC_40 TSMC_8 VDDI pch_svt_mac l=20n nfin=3 
+ m=1 
MP29<0> TSMC_41 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP29<1> TSMC_42 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP29<2> TSMC_43 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP29<3> TSMC_44 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP29<4> TSMC_45 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP29<5> TSMC_46 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP29<6> TSMC_47 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP29<7> TSMC_48 TSMC_23 VDDAI VDDI pch_svt_mac l=20n nfin=2 m=1 
XPRECHARGE<0> TSMC_1 TSMC_9 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
XPRECHARGE<1> TSMC_2 TSMC_10 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
XPRECHARGE<2> TSMC_3 TSMC_11 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
XPRECHARGE<3> TSMC_4 TSMC_12 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
XPRECHARGE<4> TSMC_5 TSMC_13 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
XPRECHARGE<5> TSMC_6 TSMC_14 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
XPRECHARGE<6> TSMC_7 TSMC_15 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
XPRECHARGE<7> TSMC_8 TSMC_16 TSMC_18 VDDI VDDI 
+ S1ALLSVTSW2000X20_PRECHARGE_M8 
MINV0_M0 TSMC_18 TSMC_17 VSSI VSSI nch_svt_mac l=20n nfin=8 m=1 
MN31_MIXV_WAS<0> TSMC_1 TSMC_49 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN31_MIXV_WAS<1> TSMC_2 TSMC_50 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN31_MIXV_WAS<2> TSMC_3 TSMC_51 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN31_MIXV_WAS<3> TSMC_4 TSMC_52 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN31_MIXV_WAS<4> TSMC_5 TSMC_53 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN31_MIXV_WAS<5> TSMC_6 TSMC_54 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN31_MIXV_WAS<6> TSMC_7 TSMC_55 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN31_MIXV_WAS<7> TSMC_8 TSMC_56 TSMC_24 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<0> TSMC_9 TSMC_49 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<1> TSMC_10 TSMC_50 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<2> TSMC_11 TSMC_51 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<3> TSMC_12 TSMC_52 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<4> TSMC_13 TSMC_53 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<5> TSMC_14 TSMC_54 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<6> TSMC_15 TSMC_55 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN18_MIXV_WAS<7> TSMC_16 TSMC_56 TSMC_22 VSSI nch_ulvt_mac l=20n nfin=5 
+ m=2 
MN13<0> TSMC_57 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN13<1> TSMC_58 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN13<2> TSMC_59 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN13<3> TSMC_60 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN13<4> TSMC_61 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN13<5> TSMC_62 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN13<6> TSMC_63 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN13<7> TSMC_64 TSMC_21 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<0> TSMC_65 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<1> TSMC_66 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<2> TSMC_67 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<3> TSMC_68 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<4> TSMC_69 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<5> TSMC_70 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<6> TSMC_71 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
MN1<7> TSMC_72 TSMC_23 VSSI VSSI nch_svt_mac l=20n nfin=3 m=1 
XI247<0> VSSI VSSI TSMC_41 TSMC_49 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI247<1> VSSI VSSI TSMC_42 TSMC_50 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI247<2> VSSI VSSI TSMC_43 TSMC_51 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI247<3> VSSI VSSI TSMC_44 TSMC_52 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI247<4> VSSI VSSI TSMC_45 TSMC_53 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI247<5> VSSI VSSI TSMC_46 TSMC_54 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI247<6> VSSI VSSI TSMC_47 TSMC_55 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI247<7> VSSI VSSI TSMC_48 TSMC_56 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=2 n_nfin=2 n_l=20n p_totalM=2 
+ p_nfin=2 p_l=20n 
XI244<0> TSMC_57 VSSI TSMC_25 TSMC_33 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI244<1> TSMC_58 VSSI TSMC_26 TSMC_34 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI244<2> TSMC_59 VSSI TSMC_27 TSMC_35 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI244<3> TSMC_60 VSSI TSMC_28 TSMC_36 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI244<4> TSMC_61 VSSI TSMC_29 TSMC_37 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI244<5> TSMC_62 VSSI TSMC_30 TSMC_38 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI244<6> TSMC_63 VSSI TSMC_31 TSMC_39 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI244<7> TSMC_64 VSSI TSMC_32 TSMC_40 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<0> TSMC_65 VSSI TSMC_25 TSMC_41 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<1> TSMC_66 VSSI TSMC_26 TSMC_42 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<2> TSMC_67 VSSI TSMC_27 TSMC_43 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<3> TSMC_68 VSSI TSMC_28 TSMC_44 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<4> TSMC_69 VSSI TSMC_29 TSMC_45 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<5> TSMC_70 VSSI TSMC_30 TSMC_46 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<6> TSMC_71 VSSI TSMC_31 TSMC_47 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI245<7> TSMC_72 VSSI TSMC_32 TSMC_48 VDDAI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    LIO_M8_NOSD
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_LIO_M8_NOSD TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 VDDAI VDDI VSSI TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
*.PININFO  TSMC_17:I TSMC_18:I TSMC_37:I TSMC_38:I TSMC_39:I TSMC_40:I 
*.PININFO  TSMC_41:I TSMC_42:I 
*.PININFO  TSMC_43:I TSMC_44:I TSMC_45:I TSMC_46:I TSMC_47:I TSMC_48:I 
*.PININFO  TSMC_49:I TSMC_50:I TSMC_51:I TSMC_52:I TSMC_53:I TSMC_54:I 
*.PININFO  TSMC_55:I TSMC_56:I TSMC_57:I TSMC_58:I TSMC_59:I TSMC_1:B 
*.PININFO  TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B 
*.PININFO  TSMC_7:B TSMC_8:B TSMC_9:B TSMC_10:B TSMC_11:B 
*.PININFO  TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B TSMC_16:B 
*.PININFO  TSMC_19:B TSMC_20:B TSMC_21:B TSMC_22:B TSMC_23:B TSMC_24:B 
*.PININFO  TSMC_25:B TSMC_26:B TSMC_27:B TSMC_28:B TSMC_29:B TSMC_30:B 
*.PININFO  TSMC_31:B TSMC_32:B TSMC_33:B TSMC_34:B TSMC_35:B TSMC_36:B VDDAI:B 
*.PININFO  VDDI:B VSSI:B 
XYPASS_U TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_18 TSMC_60 TSMC_61 TSMC_62 TSMC_63 VDDAI VDDI VSSI 
+ TSMC_64 TSMC_65 TSMC_66 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 S1ALLSVTSW2000X20_YPASS_M8_NOSD 
XYPASS_D TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_17 TSMC_67 TSMC_68 TSMC_69 TSMC_63 VDDAI VDDI VSSI TSMC_64 
+ TSMC_65 TSMC_66 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 S1ALLSVTSW2000X20_YPASS_M8_NOSD 
XIO_RWBLK TSMC_67 TSMC_60 TSMC_17 TSMC_18 TSMC_69 TSMC_62 TSMC_68 TSMC_61 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_63 TSMC_40 VDDAI VDDI 
+ VSSI TSMC_64 TSMC_41 TSMC_65 TSMC_66 S1ALLSVTSW2000X20_IO_RWBLK_M8 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    LIO_M8_S
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_LIO_M8_S TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 VDDI VSSI TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
*.PININFO  TSMC_17:I TSMC_18:I TSMC_37:I TSMC_38:I TSMC_39:I TSMC_40:I 
*.PININFO  TSMC_41:I TSMC_42:I 
*.PININFO  TSMC_43:I TSMC_44:I TSMC_45:I TSMC_46:I TSMC_47:I TSMC_48:I 
*.PININFO  TSMC_49:I TSMC_50:I TSMC_51:I TSMC_52:I TSMC_53:I TSMC_54:I 
*.PININFO  TSMC_55:I TSMC_56:I TSMC_57:I TSMC_58:I TSMC_59:I TSMC_1:B 
*.PININFO  TSMC_2:B TSMC_3:B TSMC_4:B TSMC_5:B TSMC_6:B 
*.PININFO  TSMC_7:B TSMC_8:B TSMC_9:B TSMC_10:B TSMC_11:B 
*.PININFO  TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B TSMC_16:B 
*.PININFO  TSMC_19:B TSMC_20:B TSMC_21:B TSMC_22:B TSMC_23:B TSMC_24:B 
*.PININFO  TSMC_25:B TSMC_26:B TSMC_27:B TSMC_28:B TSMC_29:B TSMC_30:B 
*.PININFO  TSMC_31:B TSMC_32:B TSMC_33:B TSMC_34:B TSMC_35:B TSMC_36:B VDDI:B 
*.PININFO  VSSI:B 
XLIO TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 VDDI VDDI VSSI 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 S1ALLSVTSW2000X20_LIO_M8_NOSD 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    LCTRL_S_M8_new_BUF_S
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_LCTRL_S_M8_new_BUF_S TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 VDDAI VDDHD VDDI TSMC_75 
+ TSMC_76 VSSI TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 
+ TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 
*.PININFO  TSMC_58:I TSMC_69:I TSMC_72:I TSMC_1:O TSMC_2:O TSMC_3:O 
*.PININFO  TSMC_40:O TSMC_41:O TSMC_42:O TSMC_43:O 
*.PININFO  TSMC_44:O TSMC_45:O TSMC_46:O TSMC_47:O 
*.PININFO  TSMC_48:O TSMC_49:O TSMC_50:O TSMC_51:O 
*.PININFO  TSMC_52:O TSMC_53:O TSMC_54:O TSMC_55:O 
*.PININFO  TSMC_60:O TSMC_61:O TSMC_63:O TSMC_64:O TSMC_67:O TSMC_68:O 
*.PININFO  TSMC_70:O TSMC_71:O TSMC_73:O TSMC_74:O TSMC_75:O TSMC_76:O 
*.PININFO  TSMC_78:O TSMC_79:O TSMC_80:O TSMC_81:O TSMC_82:O 
*.PININFO  TSMC_83:O TSMC_84:O TSMC_85:O TSMC_86:O TSMC_87:O 
*.PININFO  TSMC_92:O TSMC_93:O TSMC_4:B TSMC_5:B TSMC_6:B 
*.PININFO  TSMC_7:B TSMC_8:B TSMC_9:B TSMC_10:B TSMC_11:B 
*.PININFO  TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B TSMC_16:B 
*.PININFO  TSMC_17:B TSMC_18:B TSMC_19:B TSMC_20:B TSMC_21:B 
*.PININFO  TSMC_22:B TSMC_23:B TSMC_24:B TSMC_25:B TSMC_26:B 
*.PININFO  TSMC_27:B TSMC_28:B TSMC_29:B TSMC_30:B TSMC_31:B 
*.PININFO  TSMC_32:B TSMC_33:B TSMC_34:B TSMC_35:B TSMC_36:B TSMC_37:B 
*.PININFO  TSMC_38:B TSMC_39:B TSMC_56:B TSMC_57:B TSMC_59:B 
*.PININFO  TSMC_62:B TSMC_65:B TSMC_66:B VDDAI:B VDDHD:B VDDI:B VSSI:B 
*.PININFO  TSMC_77:B TSMC_88:B 
*.PININFO  TSMC_89:B TSMC_90:B TSMC_91:B 
MVDDHD_GG_MIXV_HD VDDHD TSMC_73 VDDI VDDI pch_svt_mac l=20n nfin=10 
+ m=32 
MVDDAI_GG_MIXV_HD TSMC_94 TSMC_3 VDDI VDDI pch_svt_mac l=20n nfin=10 
+ m=32 
XI269 VSSI VSSI TSMC_95 TSMC_71 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
XI260_MIXV_DFTUUU VSSI VSSI TSMC_72 TSMC_96 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=1 n_nfin=5 n_l=20n p_totalM=1 
+ p_nfin=5 p_l=20n 
XI262_MIXV_DFTUUU VSSI VSSI TSMC_96 TSMC_73 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=2 n_nfin=5 n_l=20n p_totalM=2 
+ p_nfin=5 p_l=20n 
XI267_MIXV_DFTUUU VSSI VSSI TSMC_97 TSMC_74 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=30 n_nfin=5 n_l=20n 
+ p_totalM=30 p_nfin=5 p_l=20n 
XI271 VSSI VSSI TSMC_98 TSMC_3 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=4 n_l=20n p_totalM=1 
+ p_nfin=4 p_l=20n 
XI265_MIXV_DFTUUU VSSI VSSI TSMC_73 TSMC_97 VDDI VDDI 
+ S1ALLSVTSW2000X20_inv_ulvt_mac_pcell_1 n_totalM=2 n_nfin=5 n_l=20n p_totalM=2 
+ p_nfin=5 p_l=20n 
XXDRV_WLP_DN TSMC_1 TSMC_99 TSMC_24 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_3 TSMC_72 TSMC_94 VDDHD VDDI VSSI TSMC_80 TSMC_81 TSMC_82 
+ TSMC_83 TSMC_88 S1ALLSVTSW2000X20_XDRV_WLP_S_M8 
XXDRV_WLP_UP TSMC_2 TSMC_100 TSMC_25 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_3 TSMC_72 TSMC_94 VDDHD VDDI VSSI TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 S1ALLSVTSW2000X20_XDRV_WLP_S_M8 
XLCTRL_BUF TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 VDDAI VDDI 
+ TSMC_75 TSMC_76 VSSI S1ALLSVTSW2000X20_LCTRL_BUF_S 
XI279 TSMC_61 TSMC_63 TSMC_76 VSSI VSSI VDDI VDDI TSMC_98 
+ S1ALLSVTSW2000X20_nor3_svt_mac_pcell_4 n_totalM=1 n_nfin=6 n_l=20n p_totalM=1 
+ p_nfin=6 p_l=20n 
XLCTRL TSMC_99 TSMC_100 TSMC_24 TSMC_25 TSMC_32 TSMC_33 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 
+ TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_72 TSMC_66 TSMC_67 TSMC_68 VDDHD 
+ VDDI VSSI TSMC_77 TSMC_78 TSMC_79 TSMC_88 TSMC_90 TSMC_91 TSMC_92 
+ TSMC_93 S1ALLSVTSW2000X20_LCTRL_M8 
XLCTRL_PM TSMC_76 TSMC_63 TSMC_64 TSMC_76 TSMC_69 TSMC_70 VDDI VSSI 
+ S1ALLSVTSW2000X20_LCTRL_PM_S 
XI258 TSMC_61 TSMC_70 VSSI VSSI VDDI VDDI TSMC_95 
+ S1ALLSVTSW2000X20_nor2_svt_mac_pcell_3 n_totalM=1 n_nfin=2 n_l=20n p_totalM=1 
+ p_nfin=2 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    LCTRL_M8_S
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_LCTRL_M8_S TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 VDDAI VDDHD VDDI TSMC_75 TSMC_76 VSSI TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 
*.PININFO  TSMC_58:I TSMC_69:I TSMC_72:I TSMC_1:O TSMC_2:O TSMC_3:O 
*.PININFO  TSMC_40:O TSMC_41:O TSMC_42:O TSMC_43:O 
*.PININFO  TSMC_44:O TSMC_45:O TSMC_46:O TSMC_47:O 
*.PININFO  TSMC_48:O TSMC_49:O TSMC_50:O TSMC_51:O 
*.PININFO  TSMC_52:O TSMC_53:O TSMC_54:O TSMC_55:O 
*.PININFO  TSMC_60:O TSMC_61:O TSMC_63:O TSMC_64:O TSMC_67:O TSMC_68:O 
*.PININFO  TSMC_70:O TSMC_71:O TSMC_73:O TSMC_74:O TSMC_75:O TSMC_76:O 
*.PININFO  TSMC_78:O TSMC_79:O TSMC_80:O TSMC_81:O TSMC_82:O 
*.PININFO  TSMC_83:O TSMC_84:O TSMC_85:O TSMC_86:O TSMC_4:B 
*.PININFO  TSMC_5:B TSMC_6:B TSMC_7:B TSMC_8:B TSMC_9:B 
*.PININFO  TSMC_10:B TSMC_11:B TSMC_12:B TSMC_13:B TSMC_14:B 
*.PININFO  TSMC_15:B TSMC_16:B TSMC_17:B TSMC_18:B TSMC_19:B 
*.PININFO  TSMC_20:B TSMC_21:B TSMC_22:B TSMC_23:B TSMC_24:B 
*.PININFO  TSMC_25:B TSMC_26:B TSMC_27:B TSMC_28:B TSMC_29:B 
*.PININFO  TSMC_30:B TSMC_31:B TSMC_32:B TSMC_33:B TSMC_34:B TSMC_35:B 
*.PININFO  TSMC_36:B TSMC_37:B TSMC_38:B TSMC_39:B TSMC_56:B 
*.PININFO  TSMC_57:B TSMC_59:B TSMC_62:B TSMC_65:B TSMC_66:B VDDAI:B VDDHD:B 
*.PININFO  VDDI:B VSSI:B TSMC_77:B TSMC_87:B TSMC_88:B 
XI257 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 
+ TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 
+ TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 
+ TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 
+ TSMC_73 TSMC_74 VDDAI VDDHD VDDI TSMC_75 TSMC_76 VSSI TSMC_77 TSMC_78 
+ TSMC_89 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 
+ TSMC_86 TSMC_87 TSMC_88 TSMC_75 TSMC_76 TSMC_90 TSMC_91 
+ S1ALLSVTSW2000X20_LCTRL_S_M8_new_BUF_S 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_LA512_SHA_NMOS
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_LA512_SHA_NMOS TSMC_1 TSMC_2 VSSI 
*.PININFO  TSMC_1:B TSMC_2:B VSSI:B 
MN5 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=2 m=4 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_LA512_SHA_A
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_LA512_SHA_A TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 VDDHD VDDI 
+ VSSI TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
*.PININFO  TSMC_37:I TSMC_40:I TSMC_45:I TSMC_46:I TSMC_47:I TSMC_43:O 
*.PININFO  TSMC_44:O TSMC_1:B TSMC_2:B TSMC_3:B TSMC_4:B 
*.PININFO  TSMC_5:B TSMC_6:B TSMC_7:B TSMC_8:B TSMC_9:B 
*.PININFO  TSMC_10:B TSMC_11:B TSMC_12:B TSMC_13:B TSMC_14:B 
*.PININFO  TSMC_15:B TSMC_16:B TSMC_17:B TSMC_18:B TSMC_19:B 
*.PININFO  TSMC_20:B TSMC_21:B TSMC_22:B TSMC_23:B TSMC_24:B 
*.PININFO  TSMC_25:B TSMC_26:B TSMC_27:B TSMC_28:B TSMC_29:B 
*.PININFO  TSMC_30:B TSMC_31:B TSMC_32:B TSMC_33:B TSMC_34:B TSMC_35:B 
*.PININFO  TSMC_36:B TSMC_38:B TSMC_39:B TSMC_41:B VDDHD:B VDDI:B VSSI:B 
*.PININFO  TSMC_42:B 
*.PININFO  TSMC_48:B TSMC_49:B TSMC_50:B 
MN7 TSMC_51 TSMC_2 TSMC_39 VSSI nch_svt_mac l=20n nfin=2 m=1 
MP9 TSMC_52 TSMC_1 TSMC_39 VSSI nch_svt_mac l=20n nfin=2 m=1 
MN0 TSMC_53 TSMC_54 TSMC_46 VSSI nch_svt_mac l=20n nfin=9 m=3 
MN6 TSMC_43 TSMC_53 VSSI VSSI nch_svt_mac l=20n nfin=10 m=8 
MM2 TSMC_44 TSMC_55 VSSI VSSI nch_svt_mac l=20n nfin=10 m=8 
MM4 TSMC_55 TSMC_56 TSMC_46 VSSI nch_svt_mac l=20n nfin=9 m=3 
MM8_MIXV_LS_UUL TSMC_53 TSMC_54 VDDI VDDI pch_lvt_mac l=20n nfin=4 m=2 
MVDDHD_GG_MIXV_HD VDDHD TSMC_40 VDDI VDDI pch_svt_mac l=20n nfin=5 m=6 
MP7 TSMC_52 TSMC_9 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MP14 TSMC_51 TSMC_2 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MM3_MIXV_LS_UUL VDDI TSMC_45 TSMC_55 VDDI pch_lvt_mac l=20n nfin=4 m=2 
MP20_MIXV_WLDV TSMC_43 TSMC_53 VDDHD VDDI pch_svt_mac l=20n nfin=18 m=8 
MP19_MIXV_LS_UUL VDDI TSMC_45 TSMC_53 VDDI pch_lvt_mac l=20n nfin=4 m=2 
MM5_MIXV_LS_UUL TSMC_55 TSMC_56 VDDI VDDI pch_lvt_mac l=20n nfin=4 m=2 
MP13 TSMC_51 TSMC_9 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
MM1_MIXV_WLDV TSMC_44 TSMC_55 VDDHD VDDI pch_svt_mac l=20n nfin=18 m=8 
MP6 TSMC_52 TSMC_1 VDDI VDDI pch_svt_mac l=20n nfin=2 m=1 
XI426 VSSI VSSI TSMC_51 TSMC_56 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
XI425 VSSI VSSI TSMC_52 TSMC_54 VDDHD VDDI 
+ S1ALLSVTSW2000X20_inv_svt_mac_pcell_1 n_totalM=1 n_nfin=3 n_l=20n p_totalM=1 
+ p_nfin=3 p_l=20n 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    XDRV_LA512_SHA_NMOS_WLPYB
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_XDRV_LA512_SHA_NMOS_WLPYB VSSI TSMC_1 TSMC_2 
*.PININFO  TSMC_1:I VSSI:B TSMC_2:B 
MN1 TSMC_2 TSMC_1 VSSI VSSI nch_svt_mac l=20n nfin=6 m=6 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WLDV_4X1_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WLDV_4X1_BASE TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 VDDHD VDDI 
+ VSSI TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I TSMC_26:I 
*.PININFO  TSMC_30:I TSMC_31:I TSMC_38:I TSMC_34:O TSMC_35:O TSMC_36:O 
*.PININFO  TSMC_37:O 
*.PININFO  TSMC_6:B TSMC_7:B TSMC_8:B TSMC_9:B TSMC_10:B 
*.PININFO  TSMC_11:B TSMC_12:B TSMC_13:B TSMC_14:B TSMC_15:B 
*.PININFO  TSMC_16:B TSMC_17:B TSMC_18:B TSMC_19:B TSMC_20:B TSMC_21:B 
*.PININFO  TSMC_22:B TSMC_23:B TSMC_24:B TSMC_25:B TSMC_27:B TSMC_28:B 
*.PININFO  TSMC_29:B 
*.PININFO  TSMC_32:B VDDHD:B VDDI:B VSSI:B TSMC_33:B TSMC_39:B TSMC_40:B 
XSHARE TSMC_5 TSMC_41 VSSI S1ALLSVTSW2000X20_XDRV_LA512_SHA_NMOS 
XWLDV_0 TSMC_1 TSMC_2 TSMC_42 TSMC_42 TSMC_42 TSMC_42 TSMC_42 TSMC_42 TSMC_5 
+ TSMC_43 TSMC_43 TSMC_43 TSMC_43 TSMC_43 TSMC_43 TSMC_43 TSMC_44 
+ TSMC_44 TSMC_44 TSMC_44 TSMC_45 TSMC_45 TSMC_45 TSMC_45 TSMC_45 
+ TSMC_45 TSMC_45 TSMC_45 TSMC_46 TSMC_46 TSMC_46 TSMC_46 TSMC_46 
+ TSMC_46 TSMC_46 TSMC_46 TSMC_26 TSMC_47 TSMC_41 TSMC_31 TSMC_48 VDDHD VDDI 
+ VSSI TSMC_49 TSMC_34 TSMC_35 TSMC_38 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_53 S1ALLSVTSW2000X20_XDRV_LA512_SHA_A 
XWLDV_1 TSMC_3 TSMC_4 TSMC_54 TSMC_54 TSMC_54 TSMC_54 TSMC_54 TSMC_54 TSMC_5 
+ TSMC_55 TSMC_55 TSMC_55 TSMC_55 TSMC_55 TSMC_55 TSMC_55 TSMC_56 
+ TSMC_56 TSMC_56 TSMC_56 TSMC_57 TSMC_57 TSMC_57 TSMC_57 TSMC_57 
+ TSMC_57 TSMC_57 TSMC_57 TSMC_58 TSMC_58 TSMC_58 TSMC_58 TSMC_58 
+ TSMC_58 TSMC_58 TSMC_58 TSMC_26 TSMC_59 TSMC_41 TSMC_31 TSMC_60 VDDHD VDDI 
+ VSSI TSMC_61 TSMC_36 TSMC_37 TSMC_38 TSMC_50 TSMC_62 TSMC_63 TSMC_64 
+ TSMC_64 S1ALLSVTSW2000X20_XDRV_LA512_SHA_A 
XI11 VSSI TSMC_38 TSMC_50 S1ALLSVTSW2000X20_XDRV_LA512_SHA_NMOS_WLPYB 
.ENDS

************************************************************************
* Library Name: N16_FFC_CHAR_MB_BOS
* Cell Name:    WLDV_4X1
* View Name:    schematic
************************************************************************

.SUBCKT S1ALLSVTSW2000X20_WLDV_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 VDDHD VDDI VSSI TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
*.PININFO  TSMC_1:I TSMC_2:I TSMC_3:I TSMC_4:I TSMC_5:I 
*.PININFO  TSMC_6:I TSMC_7:I TSMC_8:I TSMC_9:I TSMC_10:I 
*.PININFO  TSMC_11:I TSMC_12:I TSMC_13:I TSMC_14:I TSMC_15:I 
*.PININFO  TSMC_16:I TSMC_37:I TSMC_42:I TSMC_43:I TSMC_52:I 
*.PININFO  TSMC_53:I TSMC_54:I TSMC_55:I TSMC_48:O TSMC_49:O TSMC_50:O 
*.PININFO  TSMC_51:O 
*.PININFO  TSMC_17:B TSMC_18:B TSMC_19:B TSMC_20:B TSMC_21:B 
*.PININFO  TSMC_22:B TSMC_23:B TSMC_24:B TSMC_25:B TSMC_26:B 
*.PININFO  TSMC_27:B TSMC_28:B TSMC_29:B TSMC_30:B TSMC_31:B TSMC_32:B 
*.PININFO  TSMC_33:B TSMC_34:B TSMC_35:B TSMC_36:B TSMC_38:B TSMC_39:B 
*.PININFO  TSMC_40:B 
*.PININFO  TSMC_41:B TSMC_44:B TSMC_45:B TSMC_46:B VDDHD:B VDDI:B VSSI:B 
*.PININFO  TSMC_47:B 
*.PININFO  TSMC_56:B TSMC_57:B TSMC_58:B TSMC_59:B 
XWLDV_4X1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_9 TSMC_17 TSMC_18 TSMC_19 
+ TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 TSMC_27 
+ TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_42 TSMC_43 TSMC_46 VDDHD 
+ VDDI VSSI TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_56 
+ TSMC_57 S1ALLSVTSW2000X20_WLDV_4X1_BASE 
.ENDS




**** End of leaf cells

.SUBCKT S1ALLSVTSW2000X20_CELL_ARR_Y TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_21 TSMC_22 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 
+ TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 
+ TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 
+ TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 
+ TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 
XMCB_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_21 TSMC_22 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_1 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_23 TSMC_24 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_25 TSMC_26 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_3 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_27 TSMC_28 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_29 TSMC_30 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_5 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_31 TSMC_32 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_33 TSMC_34 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_7 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_35 TSMC_36 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_37 TSMC_38 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_9 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_39 TSMC_40 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_10 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_41 TSMC_42 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_11 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_43 TSMC_44 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_12 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_45 TSMC_46 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_13 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_47 TSMC_48 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_14 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_49 TSMC_50 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_15 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_51 TSMC_52 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_16 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_53 TSMC_54 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_17 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_55 TSMC_56 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_18 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_57 TSMC_58 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_19 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_59 TSMC_60 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_20 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_61 TSMC_62 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_21 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_63 TSMC_64 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_22 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_65 TSMC_66 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_23 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_67 TSMC_68 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_24 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_69 TSMC_70 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_25 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_71 TSMC_72 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_26 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_73 TSMC_74 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_27 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_75 TSMC_76 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_28 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_77 TSMC_78 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_29 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_79 TSMC_80 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_30 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_81 TSMC_82 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_31 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_83 TSMC_84 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_32 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_85 TSMC_86 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_33 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_87 TSMC_88 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_34 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_89 TSMC_90 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_35 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_91 TSMC_92 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_36 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_93 TSMC_94 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_37 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_95 TSMC_96 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_38 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_97 TSMC_98 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_39 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_99 TSMC_100 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_40 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_101 TSMC_102 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_41 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_103 TSMC_104 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_42 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_105 TSMC_106 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_43 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_107 TSMC_108 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_44 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_109 TSMC_110 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_45 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_111 TSMC_112 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_46 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_113 TSMC_114 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_47 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_115 TSMC_116 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_48 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_117 TSMC_118 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_49 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_119 TSMC_120 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_50 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_121 TSMC_122 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_51 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_123 TSMC_124 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_52 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_125 TSMC_126 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_53 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_127 TSMC_128 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_54 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_129 TSMC_130 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_55 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_131 TSMC_132 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_56 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_133 TSMC_134 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_57 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_135 TSMC_136 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_58 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_137 TSMC_138 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_59 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_139 TSMC_140 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_60 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_141 TSMC_142 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_61 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_143 TSMC_144 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_62 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_145 TSMC_146 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_63 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_147 TSMC_148 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_64 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_149 TSMC_150 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_65 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_151 TSMC_152 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_66 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_153 TSMC_154 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_67 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_155 TSMC_156 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_68 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_157 TSMC_158 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_69 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_159 TSMC_160 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_70 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_161 TSMC_162 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_71 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_163 TSMC_164 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_72 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_165 TSMC_166 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_73 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_167 TSMC_168 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_74 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_169 TSMC_170 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_75 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_171 TSMC_172 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_76 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_173 TSMC_174 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_77 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_175 TSMC_176 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_78 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_177 TSMC_178 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_79 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_179 TSMC_180 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_80 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_181 TSMC_182 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_81 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_183 TSMC_184 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_82 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_185 TSMC_186 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_83 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_187 TSMC_188 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_84 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_189 TSMC_190 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_85 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_191 TSMC_192 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_86 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_193 TSMC_194 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_87 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_195 TSMC_196 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_88 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_197 TSMC_198 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_89 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_199 TSMC_200 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_90 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_201 TSMC_202 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_91 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_203 TSMC_204 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_92 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_205 TSMC_206 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_93 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_207 TSMC_208 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_94 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_209 TSMC_210 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_95 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_211 TSMC_212 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_96 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_213 TSMC_214 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_97 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_215 TSMC_216 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_98 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_217 TSMC_218 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_99 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_219 TSMC_220 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_100 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_221 TSMC_222 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_101 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_223 TSMC_224 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_102 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_225 TSMC_226 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_103 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_227 TSMC_228 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_104 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_229 TSMC_230 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_105 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_231 TSMC_232 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_106 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_233 TSMC_234 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_107 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_235 TSMC_236 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_108 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_237 TSMC_238 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_109 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_239 TSMC_240 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_110 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_241 TSMC_242 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_111 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_243 TSMC_244 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_112 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_245 TSMC_246 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_113 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_247 TSMC_248 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_114 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_249 TSMC_250 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_115 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_251 TSMC_252 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_116 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_253 TSMC_254 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_117 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_255 TSMC_256 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_118 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_257 TSMC_258 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_119 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_259 TSMC_260 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_120 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_261 TSMC_262 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_121 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_263 TSMC_264 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_122 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_265 TSMC_266 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_123 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_267 TSMC_268 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_124 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_269 TSMC_270 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_125 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_271 TSMC_272 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_126 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_273 TSMC_274 
+ S1ALLSVTSW2000X20_MCB_2X8 
XMCB_127 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 VDDAI VDDI VSSI TSMC_275 TSMC_276 
+ S1ALLSVTSW2000X20_MCB_2X8 
.ENDS

.SUBCKT S1ALLSVTSW2000X20_WLDV_F_DN TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 VDDHD VDDI VSSI TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 
+ TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 
+ TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 
+ TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 
+ TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 
+ TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 
+ TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
XWLDV_4X1_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_1 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_3 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_5 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_7 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_9 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_10 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_11 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_12 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_13 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_14 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_15 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_16 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_17 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_18 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_19 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_20 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_21 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_22 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_23 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_24 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_25 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_26 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_27 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_28 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_29 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_30 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_31 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_32 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_33 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_34 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_35 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_36 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_37 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_38 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_39 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_40 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_41 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_42 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_43 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_44 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_45 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_46 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_47 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_48 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_49 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_50 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_51 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_52 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_53 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_54 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_55 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_56 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_57 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_58 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_59 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_60 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_61 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_62 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_294 TSMC_295 TSMC_296 TSMC_297 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_63 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
.ENDS

.SUBCKT S1ALLSVTSW2000X20_WLDV_F TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 VDDHD VDDI VSSI TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 
+ TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 
+ TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 
+ TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 
+ TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 
+ TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 
+ TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 
+ TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 
+ TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 
+ TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 
+ TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 
+ TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 
+ TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 
+ TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 
+ TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 
+ TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 
+ TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 
+ TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 
+ TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 
+ TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 
+ TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
XWLDV_4X1_0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_1 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_2 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_3 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_4 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_5 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_6 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_7 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_9 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_10 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_11 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_12 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_13 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_302 TSMC_303 TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_14 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_15 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_16 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_17 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_18 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_19 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_20 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_21 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_22 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_23 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_24 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_25 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_26 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_27 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_28 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_29 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_30 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_31 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_303 TSMC_302 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_32 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_33 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_34 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_35 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_36 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_37 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_38 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_39 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_40 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_41 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_42 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_43 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_44 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_45 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_46 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_47 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_304 TSMC_302 
+ TSMC_303 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_48 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_49 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_50 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_51 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_10 TSMC_9 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_52 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_53 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_11 TSMC_9 TSMC_10 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_54 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_55 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_12 TSMC_9 TSMC_10 TSMC_11 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_56 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_57 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_13 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_58 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_59 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_14 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_60 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_61 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_15 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_62 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_294 TSMC_295 TSMC_296 TSMC_297 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
XWLDV_4X1_63 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_1 TSMC_2 TSMC_3 TSMC_4 
+ TSMC_16 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 
+ TSMC_33 TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 
+ TSMC_41 TSMC_42 TSMC_43 TSMC_310 TSMC_311 TSMC_44 VDDHD VDDI VSSI 
+ TSMC_45 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_305 TSMC_302 
+ TSMC_303 TSMC_304 TSMC_306 TSMC_307 TSMC_308 TSMC_309 
+ S1ALLSVTSW2000X20_WLDV_4X1 
.ENDS

.SUBCKT S1ALLSVTSW2000X20_GTRK_ARR TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 VDDAI VDDI VSSI TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 
+ TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 
+ TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 
+ TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 
+ TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 
+ TSMC_168 TSMC_169 TSMC_170 TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 
+ TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 
+ TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 
+ TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 
+ TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 
+ TSMC_232 TSMC_233 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 
+ TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 
+ TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 
+ TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 
+ TSMC_296 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
+ TSMC_312 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 
+ TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 
+ TSMC_328 TSMC_329 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 
+ TSMC_336 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 
+ TSMC_344 TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 
+ TSMC_352 TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 
+ TSMC_360 TSMC_361 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 
+ TSMC_384 TSMC_385 TSMC_386 TSMC_387 
XTRKBL_OFF_127 TSMC_129 VDDI VDDAI VSSI TSMC_131 TSMC_132 TSMC_388 
+ TSMC_389 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_126 TSMC_129 VDDI VDDAI VSSI TSMC_133 TSMC_134 TSMC_390 
+ TSMC_388 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_125 TSMC_129 VDDI VDDAI VSSI TSMC_135 TSMC_136 TSMC_391 
+ TSMC_390 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_124 TSMC_129 VDDI VDDAI VSSI TSMC_137 TSMC_138 TSMC_392 
+ TSMC_391 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_123 TSMC_129 VDDI VDDAI VSSI TSMC_139 TSMC_140 TSMC_393 
+ TSMC_392 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_122 TSMC_129 VDDI VDDAI VSSI TSMC_141 TSMC_142 TSMC_394 
+ TSMC_393 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_121 TSMC_129 VDDI VDDAI VSSI TSMC_143 TSMC_144 TSMC_395 
+ TSMC_394 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_120 TSMC_129 VDDI VDDAI VSSI TSMC_145 TSMC_146 TSMC_396 
+ TSMC_395 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_119 TSMC_129 VDDI VDDAI VSSI TSMC_147 TSMC_148 TSMC_397 
+ TSMC_396 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_118 TSMC_129 VDDI VDDAI VSSI TSMC_149 TSMC_150 TSMC_398 
+ TSMC_397 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_117 TSMC_129 VDDI VDDAI VSSI TSMC_151 TSMC_152 TSMC_399 
+ TSMC_398 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_116 TSMC_129 VDDI VDDAI VSSI TSMC_153 TSMC_154 TSMC_400 
+ TSMC_399 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_115 TSMC_129 VDDI VDDAI VSSI TSMC_155 TSMC_156 TSMC_401 
+ TSMC_400 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_114 TSMC_129 VDDI VDDAI VSSI TSMC_157 TSMC_158 TSMC_402 
+ TSMC_401 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_113 TSMC_129 VDDI VDDAI VSSI TSMC_159 TSMC_160 TSMC_403 
+ TSMC_402 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_112 TSMC_129 VDDI VDDAI VSSI TSMC_161 TSMC_162 TSMC_404 
+ TSMC_403 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_111 TSMC_129 VDDI VDDAI VSSI TSMC_163 TSMC_164 TSMC_405 
+ TSMC_404 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_110 TSMC_129 VDDI VDDAI VSSI TSMC_165 TSMC_166 TSMC_406 
+ TSMC_405 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_109 TSMC_129 VDDI VDDAI VSSI TSMC_167 TSMC_168 TSMC_407 
+ TSMC_406 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_108 TSMC_129 VDDI VDDAI VSSI TSMC_169 TSMC_170 TSMC_408 
+ TSMC_407 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_107 TSMC_129 VDDI VDDAI VSSI TSMC_171 TSMC_172 TSMC_409 
+ TSMC_408 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_106 TSMC_129 VDDI VDDAI VSSI TSMC_173 TSMC_174 TSMC_410 
+ TSMC_409 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_105 TSMC_129 VDDI VDDAI VSSI TSMC_175 TSMC_176 TSMC_411 
+ TSMC_410 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_104 TSMC_129 VDDI VDDAI VSSI TSMC_177 TSMC_178 TSMC_412 
+ TSMC_411 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_103 TSMC_129 VDDI VDDAI VSSI TSMC_179 TSMC_180 TSMC_413 
+ TSMC_412 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_102 TSMC_129 VDDI VDDAI VSSI TSMC_181 TSMC_182 TSMC_414 
+ TSMC_413 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_101 TSMC_129 VDDI VDDAI VSSI TSMC_183 TSMC_184 TSMC_415 
+ TSMC_414 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_100 TSMC_129 VDDI VDDAI VSSI TSMC_185 TSMC_186 TSMC_416 
+ TSMC_415 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_99 TSMC_129 VDDI VDDAI VSSI TSMC_187 TSMC_188 TSMC_417 
+ TSMC_416 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_98 TSMC_129 VDDI VDDAI VSSI TSMC_189 TSMC_190 TSMC_418 
+ TSMC_417 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_97 TSMC_129 VDDI VDDAI VSSI TSMC_191 TSMC_192 TSMC_419 
+ TSMC_418 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_96 TSMC_129 VDDI VDDAI VSSI TSMC_193 TSMC_194 TSMC_420 
+ TSMC_419 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_95 TSMC_129 VDDI VDDAI VSSI TSMC_195 TSMC_196 TSMC_421 
+ TSMC_420 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_94 TSMC_129 VDDI VDDAI VSSI TSMC_197 TSMC_198 TSMC_422 
+ TSMC_421 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_93 TSMC_129 VDDI VDDAI VSSI TSMC_199 TSMC_200 TSMC_423 
+ TSMC_422 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_92 TSMC_129 VDDI VDDAI VSSI TSMC_201 TSMC_202 TSMC_424 
+ TSMC_423 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_91 TSMC_129 VDDI VDDAI VSSI TSMC_203 TSMC_204 TSMC_425 
+ TSMC_424 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_90 TSMC_129 VDDI VDDAI VSSI TSMC_205 TSMC_206 TSMC_426 
+ TSMC_425 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_89 TSMC_129 VDDI VDDAI VSSI TSMC_207 TSMC_208 TSMC_427 
+ TSMC_426 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_88 TSMC_129 VDDI VDDAI VSSI TSMC_209 TSMC_210 TSMC_428 
+ TSMC_427 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_87 TSMC_129 VDDI VDDAI VSSI TSMC_211 TSMC_212 TSMC_429 
+ TSMC_428 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_86 TSMC_129 VDDI VDDAI VSSI TSMC_213 TSMC_214 TSMC_430 
+ TSMC_429 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_85 TSMC_129 VDDI VDDAI VSSI TSMC_215 TSMC_216 TSMC_431 
+ TSMC_430 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_84 TSMC_129 VDDI VDDAI VSSI TSMC_217 TSMC_218 TSMC_432 
+ TSMC_431 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_83 TSMC_129 VDDI VDDAI VSSI TSMC_219 TSMC_220 TSMC_433 
+ TSMC_432 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_82 TSMC_129 VDDI VDDAI VSSI TSMC_221 TSMC_222 TSMC_434 
+ TSMC_433 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_81 TSMC_129 VDDI VDDAI VSSI TSMC_223 TSMC_224 TSMC_435 
+ TSMC_434 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_80 TSMC_129 VDDI VDDAI VSSI TSMC_225 TSMC_226 TSMC_436 
+ TSMC_435 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_79 TSMC_129 VDDI VDDAI VSSI TSMC_227 TSMC_228 TSMC_437 
+ TSMC_436 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_78 TSMC_129 VDDI VDDAI VSSI TSMC_229 TSMC_230 TSMC_438 
+ TSMC_437 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_77 TSMC_129 VDDI VDDAI VSSI TSMC_231 TSMC_232 TSMC_439 
+ TSMC_438 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_76 TSMC_129 VDDI VDDAI VSSI TSMC_233 TSMC_234 TSMC_440 
+ TSMC_439 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_75 TSMC_129 VDDI VDDAI VSSI TSMC_235 TSMC_236 TSMC_441 
+ TSMC_440 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_74 TSMC_129 VDDI VDDAI VSSI TSMC_237 TSMC_238 TSMC_442 
+ TSMC_441 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_73 TSMC_129 VDDI VDDAI VSSI TSMC_239 TSMC_240 TSMC_443 
+ TSMC_442 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_72 TSMC_129 VDDI VDDAI VSSI TSMC_241 TSMC_242 TSMC_444 
+ TSMC_443 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_71 TSMC_129 VDDI VDDAI VSSI TSMC_243 TSMC_244 TSMC_445 
+ TSMC_444 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_70 TSMC_129 VDDI VDDAI VSSI TSMC_245 TSMC_246 TSMC_446 
+ TSMC_445 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_69 TSMC_129 VDDI VDDAI VSSI TSMC_247 TSMC_248 TSMC_447 
+ TSMC_446 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_68 TSMC_129 VDDI VDDAI VSSI TSMC_249 TSMC_250 TSMC_448 
+ TSMC_447 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_67 TSMC_129 VDDI VDDAI VSSI TSMC_251 TSMC_252 TSMC_449 
+ TSMC_448 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_66 TSMC_129 VDDI VDDAI VSSI TSMC_253 TSMC_254 TSMC_450 
+ TSMC_449 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_65 TSMC_129 VDDI VDDAI VSSI TSMC_255 TSMC_256 TSMC_451 
+ TSMC_450 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_64 TSMC_129 VDDI VDDAI VSSI TSMC_257 TSMC_258 TSMC_452 
+ TSMC_451 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_63 TSMC_129 VDDI VDDAI VSSI TSMC_259 TSMC_260 TSMC_453 
+ TSMC_452 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_62 TSMC_129 VDDI VDDAI VSSI TSMC_261 TSMC_262 TSMC_454 
+ TSMC_453 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_61 TSMC_129 VDDI VDDAI VSSI TSMC_263 TSMC_264 TSMC_455 
+ TSMC_454 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_60 TSMC_129 VDDI VDDAI VSSI TSMC_265 TSMC_266 TSMC_456 
+ TSMC_455 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_59 TSMC_129 VDDI VDDAI VSSI TSMC_267 TSMC_268 TSMC_457 
+ TSMC_456 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_58 TSMC_129 VDDI VDDAI VSSI TSMC_269 TSMC_270 TSMC_458 
+ TSMC_457 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_57 TSMC_129 VDDI VDDAI VSSI TSMC_271 TSMC_272 TSMC_459 
+ TSMC_458 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_56 TSMC_129 VDDI VDDAI VSSI TSMC_273 TSMC_274 TSMC_460 
+ TSMC_459 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_55 TSMC_129 VDDI VDDAI VSSI TSMC_275 TSMC_276 TSMC_461 
+ TSMC_460 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_54 TSMC_129 VDDI VDDAI VSSI TSMC_277 TSMC_278 TSMC_462 
+ TSMC_461 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_53 TSMC_129 VDDI VDDAI VSSI TSMC_279 TSMC_280 TSMC_463 
+ TSMC_462 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_52 TSMC_129 VDDI VDDAI VSSI TSMC_281 TSMC_282 TSMC_464 
+ TSMC_463 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_51 TSMC_129 VDDI VDDAI VSSI TSMC_283 TSMC_284 TSMC_465 
+ TSMC_464 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_50 TSMC_129 VDDI VDDAI VSSI TSMC_285 TSMC_286 TSMC_466 
+ TSMC_465 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_49 TSMC_129 VDDI VDDAI VSSI TSMC_287 TSMC_288 TSMC_467 
+ TSMC_466 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_48 TSMC_129 VDDI VDDAI VSSI TSMC_289 TSMC_290 TSMC_468 
+ TSMC_467 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_47 TSMC_129 VDDI VDDAI VSSI TSMC_291 TSMC_292 TSMC_469 
+ TSMC_468 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_46 TSMC_129 VDDI VDDAI VSSI TSMC_293 TSMC_294 TSMC_470 
+ TSMC_469 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_45 TSMC_129 VDDI VDDAI VSSI TSMC_295 TSMC_296 TSMC_471 
+ TSMC_470 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_44 TSMC_129 VDDI VDDAI VSSI TSMC_297 TSMC_298 TSMC_472 
+ TSMC_471 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_43 TSMC_129 VDDI VDDAI VSSI TSMC_299 TSMC_300 TSMC_473 
+ TSMC_472 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_42 TSMC_129 VDDI VDDAI VSSI TSMC_301 TSMC_302 TSMC_474 
+ TSMC_473 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_41 TSMC_129 VDDI VDDAI VSSI TSMC_303 TSMC_304 TSMC_475 
+ TSMC_474 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_40 TSMC_129 VDDI VDDAI VSSI TSMC_305 TSMC_306 TSMC_476 
+ TSMC_475 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_39 TSMC_129 VDDI VDDAI VSSI TSMC_307 TSMC_308 TSMC_477 
+ TSMC_476 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_38 TSMC_129 VDDI VDDAI VSSI TSMC_309 TSMC_310 TSMC_478 
+ TSMC_477 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_37 TSMC_129 VDDI VDDAI VSSI TSMC_311 TSMC_312 TSMC_479 
+ TSMC_478 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_36 TSMC_129 VDDI VDDAI VSSI TSMC_313 TSMC_314 TSMC_480 
+ TSMC_479 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_35 TSMC_129 VDDI VDDAI VSSI TSMC_315 TSMC_316 TSMC_481 
+ TSMC_480 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_34 TSMC_129 VDDI VDDAI VSSI TSMC_317 TSMC_318 TSMC_482 
+ TSMC_481 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_33 TSMC_129 VDDI VDDAI VSSI TSMC_319 TSMC_320 TSMC_483 
+ TSMC_482 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_32 TSMC_129 VDDI VDDAI VSSI TSMC_321 TSMC_322 TSMC_484 
+ TSMC_483 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_31 TSMC_129 VDDI VDDAI VSSI TSMC_323 TSMC_324 TSMC_485 
+ TSMC_484 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_30 TSMC_129 VDDI VDDAI VSSI TSMC_325 TSMC_326 TSMC_486 
+ TSMC_485 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_29 TSMC_129 VDDI VDDAI VSSI TSMC_327 TSMC_328 TSMC_487 
+ TSMC_486 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_28 TSMC_129 VDDI VDDAI VSSI TSMC_329 TSMC_330 TSMC_488 
+ TSMC_487 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_27 TSMC_129 VDDI VDDAI VSSI TSMC_331 TSMC_332 TSMC_489 
+ TSMC_488 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_26 TSMC_129 VDDI VDDAI VSSI TSMC_333 TSMC_334 TSMC_490 
+ TSMC_489 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_25 TSMC_129 VDDI VDDAI VSSI TSMC_335 TSMC_336 TSMC_491 
+ TSMC_490 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_24 TSMC_129 VDDI VDDAI VSSI TSMC_337 TSMC_338 TSMC_492 
+ TSMC_491 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_23 TSMC_129 VDDI VDDAI VSSI TSMC_339 TSMC_340 TSMC_493 
+ TSMC_492 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_22 TSMC_129 VDDI VDDAI VSSI TSMC_341 TSMC_342 TSMC_494 
+ TSMC_493 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_21 TSMC_129 VDDI VDDAI VSSI TSMC_343 TSMC_344 TSMC_495 
+ TSMC_494 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_20 TSMC_129 VDDI VDDAI VSSI TSMC_345 TSMC_346 TSMC_496 
+ TSMC_495 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_19 TSMC_129 VDDI VDDAI VSSI TSMC_347 TSMC_348 TSMC_497 
+ TSMC_496 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_18 TSMC_129 VDDI VDDAI VSSI TSMC_349 TSMC_350 TSMC_498 
+ TSMC_497 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_17 TSMC_129 VDDI VDDAI VSSI TSMC_351 TSMC_352 TSMC_499 
+ TSMC_498 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_OFF_16 TSMC_129 VDDI VDDAI VSSI TSMC_353 TSMC_354 TSMC_500 
+ TSMC_499 S1ALLSVTSW2000X20_TRKBL_OFF_X2 
XTRKBL_ISO_15 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_355 TSMC_356 
+ TSMC_500 S1ALLSVTSW2000X20_TRKBL_ISO_X2 
XTRKBL_ON_14 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_357 
+ TSMC_358 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_13 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_359 
+ TSMC_360 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_12 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_361 
+ TSMC_362 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_11 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_363 
+ TSMC_364 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_10 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_365 
+ TSMC_366 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_9 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_367 
+ TSMC_368 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_8 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_369 
+ TSMC_370 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_7 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_371 
+ TSMC_372 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_6 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_373 
+ TSMC_374 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_5 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_375 
+ TSMC_376 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_4 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_377 
+ TSMC_378 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_3 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_379 
+ TSMC_380 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_2 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_381 
+ TSMC_382 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_1 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_383 
+ TSMC_384 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRKBL_ON_0 TSMC_129 TSMC_387 TSMC_387 VDDI VDDAI VSSI TSMC_385 
+ TSMC_386 S1ALLSVTSW2000X20_TRKBL_ON_X2 
XTRK_PRE TSMC_130 TSMC_129 TSMC_387 VDDAI VDDI VSSI TSMC_501 TSMC_502 
+ S1ALLSVTSW2000X20_TKBL_TRKPRE 
.ENDS

.SUBCKT S1ALLSVTSW2000X20_BANK0_F TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 VDDAI VDDHD VDDI VSSI TSMC_173 TSMC_174 TSMC_175 
+ TSMC_176 TSMC_177 TSMC_178 
XLIO_M8_S_AL_0 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 
+ TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 
+ TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 TSMC_36 
+ TSMC_68 TSMC_100 TSMC_132 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_1 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 
+ TSMC_247 TSMC_248 TSMC_249 TSMC_195 TSMC_196 TSMC_250 TSMC_251 
+ TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 
+ TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_37 
+ TSMC_69 TSMC_101 TSMC_133 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_2 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 TSMC_273 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 
+ TSMC_279 TSMC_280 TSMC_281 TSMC_195 TSMC_196 TSMC_282 TSMC_283 
+ TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 
+ TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 TSMC_38 
+ TSMC_70 TSMC_102 TSMC_134 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_3 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 
+ TSMC_311 TSMC_312 TSMC_313 TSMC_195 TSMC_196 TSMC_314 TSMC_315 
+ TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 TSMC_321 TSMC_322 
+ TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_39 
+ TSMC_71 TSMC_103 TSMC_135 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_4 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 
+ TSMC_336 TSMC_337 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 
+ TSMC_343 TSMC_344 TSMC_345 TSMC_195 TSMC_196 TSMC_346 TSMC_347 
+ TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 
+ TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 TSMC_361 TSMC_40 
+ TSMC_72 TSMC_104 TSMC_136 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_5 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 
+ TSMC_375 TSMC_376 TSMC_377 TSMC_195 TSMC_196 TSMC_378 TSMC_379 
+ TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 TSMC_385 TSMC_386 
+ TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_41 
+ TSMC_73 TSMC_105 TSMC_137 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_6 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 
+ TSMC_400 TSMC_401 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 
+ TSMC_407 TSMC_408 TSMC_409 TSMC_195 TSMC_196 TSMC_410 TSMC_411 
+ TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 
+ TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 TSMC_425 TSMC_42 
+ TSMC_74 TSMC_106 TSMC_138 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_7 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 
+ TSMC_432 TSMC_433 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 
+ TSMC_439 TSMC_440 TSMC_441 TSMC_195 TSMC_196 TSMC_442 TSMC_443 
+ TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 TSMC_449 TSMC_450 
+ TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 TSMC_457 TSMC_43 
+ TSMC_75 TSMC_107 TSMC_139 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_8 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 
+ TSMC_464 TSMC_465 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 
+ TSMC_471 TSMC_472 TSMC_473 TSMC_195 TSMC_196 TSMC_474 TSMC_475 
+ TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 
+ TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 TSMC_489 TSMC_44 
+ TSMC_76 TSMC_108 TSMC_140 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_9 TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 
+ TSMC_496 TSMC_497 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 
+ TSMC_503 TSMC_504 TSMC_505 TSMC_195 TSMC_196 TSMC_506 TSMC_507 
+ TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 TSMC_513 TSMC_514 
+ TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_45 
+ TSMC_77 TSMC_109 TSMC_141 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_10 TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 TSMC_527 
+ TSMC_528 TSMC_529 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 
+ TSMC_535 TSMC_536 TSMC_537 TSMC_195 TSMC_196 TSMC_538 TSMC_539 
+ TSMC_540 TSMC_541 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 
+ TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 TSMC_552 TSMC_553 
+ TSMC_46 TSMC_78 TSMC_110 TSMC_142 TSMC_213 TSMC_214 VDDI VSSI 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_ABL_11 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 TSMC_559 
+ TSMC_560 TSMC_561 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_195 TSMC_196 TSMC_570 TSMC_571 
+ TSMC_572 TSMC_573 TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 
+ TSMC_579 TSMC_580 TSMC_581 TSMC_582 TSMC_583 TSMC_584 TSMC_585 
+ TSMC_47 TSMC_79 TSMC_111 TSMC_143 TSMC_213 TSMC_214 VDDI VSSI 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CL_12 TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 TSMC_591 
+ TSMC_592 TSMC_593 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 TSMC_601 TSMC_195 TSMC_196 TSMC_602 TSMC_603 
+ TSMC_604 TSMC_605 TSMC_606 TSMC_607 TSMC_608 TSMC_609 TSMC_610 
+ TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 TSMC_616 TSMC_617 
+ TSMC_48 TSMC_80 TSMC_112 TSMC_144 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CL_13 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 TSMC_623 
+ TSMC_624 TSMC_625 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 TSMC_633 TSMC_195 TSMC_196 TSMC_634 TSMC_635 
+ TSMC_636 TSMC_637 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 
+ TSMC_643 TSMC_644 TSMC_645 TSMC_646 TSMC_647 TSMC_648 TSMC_649 
+ TSMC_49 TSMC_81 TSMC_113 TSMC_145 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CL_14 TSMC_650 TSMC_651 TSMC_652 TSMC_653 TSMC_654 TSMC_655 
+ TSMC_656 TSMC_657 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 
+ TSMC_663 TSMC_664 TSMC_665 TSMC_195 TSMC_196 TSMC_666 TSMC_667 
+ TSMC_668 TSMC_669 TSMC_670 TSMC_671 TSMC_672 TSMC_673 TSMC_674 
+ TSMC_675 TSMC_676 TSMC_677 TSMC_678 TSMC_679 TSMC_680 TSMC_681 
+ TSMC_50 TSMC_82 TSMC_114 TSMC_146 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CBL_L_15 TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 
+ TSMC_687 TSMC_688 TSMC_689 TSMC_690 TSMC_691 TSMC_692 TSMC_693 
+ TSMC_694 TSMC_695 TSMC_696 TSMC_697 TSMC_195 TSMC_196 TSMC_698 
+ TSMC_699 TSMC_700 TSMC_701 TSMC_702 TSMC_703 TSMC_704 TSMC_705 
+ TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 TSMC_711 TSMC_712 
+ TSMC_713 TSMC_51 TSMC_83 TSMC_115 TSMC_147 TSMC_213 TSMC_214 VDDI VSSI 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CBL_R_16 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 
+ TSMC_719 TSMC_720 TSMC_721 TSMC_722 TSMC_723 TSMC_724 TSMC_725 
+ TSMC_726 TSMC_727 TSMC_728 TSMC_729 TSMC_195 TSMC_196 TSMC_730 
+ TSMC_731 TSMC_732 TSMC_733 TSMC_734 TSMC_735 TSMC_736 TSMC_737 
+ TSMC_738 TSMC_739 TSMC_740 TSMC_741 TSMC_742 TSMC_743 TSMC_744 
+ TSMC_745 TSMC_52 TSMC_84 TSMC_116 TSMC_148 TSMC_213 TSMC_214 VDDI VSSI 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_C_R_17 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 TSMC_751 
+ TSMC_752 TSMC_753 TSMC_754 TSMC_755 TSMC_756 TSMC_757 TSMC_758 
+ TSMC_759 TSMC_760 TSMC_761 TSMC_195 TSMC_196 TSMC_762 TSMC_763 
+ TSMC_764 TSMC_765 TSMC_766 TSMC_767 TSMC_768 TSMC_769 TSMC_770 
+ TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_775 TSMC_776 TSMC_777 
+ TSMC_53 TSMC_85 TSMC_117 TSMC_149 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_C_R_18 TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_782 TSMC_783 
+ TSMC_784 TSMC_785 TSMC_786 TSMC_787 TSMC_788 TSMC_789 TSMC_790 
+ TSMC_791 TSMC_792 TSMC_793 TSMC_195 TSMC_196 TSMC_794 TSMC_795 
+ TSMC_796 TSMC_797 TSMC_798 TSMC_799 TSMC_800 TSMC_801 TSMC_802 
+ TSMC_803 TSMC_804 TSMC_805 TSMC_806 TSMC_807 TSMC_808 TSMC_809 
+ TSMC_54 TSMC_86 TSMC_118 TSMC_150 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_C_R_19 TSMC_810 TSMC_811 TSMC_812 TSMC_813 TSMC_814 TSMC_815 
+ TSMC_816 TSMC_817 TSMC_818 TSMC_819 TSMC_820 TSMC_821 TSMC_822 
+ TSMC_823 TSMC_824 TSMC_825 TSMC_195 TSMC_196 TSMC_826 TSMC_827 
+ TSMC_828 TSMC_829 TSMC_830 TSMC_831 TSMC_832 TSMC_833 TSMC_834 
+ TSMC_835 TSMC_836 TSMC_837 TSMC_838 TSMC_839 TSMC_840 TSMC_841 
+ TSMC_55 TSMC_87 TSMC_119 TSMC_151 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_ABL_R_20 TSMC_842 TSMC_843 TSMC_844 TSMC_845 TSMC_846 
+ TSMC_847 TSMC_848 TSMC_849 TSMC_850 TSMC_851 TSMC_852 TSMC_853 
+ TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_195 TSMC_196 TSMC_858 
+ TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 TSMC_864 TSMC_865 
+ TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 TSMC_872 
+ TSMC_873 TSMC_56 TSMC_88 TSMC_120 TSMC_152 TSMC_213 TSMC_214 VDDI VSSI 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_21 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 
+ TSMC_880 TSMC_881 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 
+ TSMC_887 TSMC_888 TSMC_889 TSMC_195 TSMC_196 TSMC_890 TSMC_891 
+ TSMC_892 TSMC_893 TSMC_894 TSMC_895 TSMC_896 TSMC_897 TSMC_898 
+ TSMC_899 TSMC_900 TSMC_901 TSMC_902 TSMC_903 TSMC_904 TSMC_905 
+ TSMC_57 TSMC_89 TSMC_121 TSMC_153 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_22 TSMC_906 TSMC_907 TSMC_908 TSMC_909 TSMC_910 TSMC_911 
+ TSMC_912 TSMC_913 TSMC_914 TSMC_915 TSMC_916 TSMC_917 TSMC_918 
+ TSMC_919 TSMC_920 TSMC_921 TSMC_195 TSMC_196 TSMC_922 TSMC_923 
+ TSMC_924 TSMC_925 TSMC_926 TSMC_927 TSMC_928 TSMC_929 TSMC_930 
+ TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 TSMC_936 TSMC_937 
+ TSMC_58 TSMC_90 TSMC_122 TSMC_154 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_23 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_195 TSMC_196 TSMC_954 TSMC_955 
+ TSMC_956 TSMC_957 TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 
+ TSMC_963 TSMC_964 TSMC_965 TSMC_966 TSMC_967 TSMC_968 TSMC_969 
+ TSMC_59 TSMC_91 TSMC_123 TSMC_155 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_24 TSMC_970 TSMC_971 TSMC_972 TSMC_973 TSMC_974 TSMC_975 
+ TSMC_976 TSMC_977 TSMC_978 TSMC_979 TSMC_980 TSMC_981 TSMC_982 
+ TSMC_983 TSMC_984 TSMC_985 TSMC_195 TSMC_196 TSMC_986 TSMC_987 
+ TSMC_988 TSMC_989 TSMC_990 TSMC_991 TSMC_992 TSMC_993 TSMC_994 
+ TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 TSMC_1000 TSMC_1001 
+ TSMC_60 TSMC_92 TSMC_124 TSMC_156 TSMC_213 TSMC_214 VDDI VSSI TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ TSMC_230 TSMC_231 TSMC_232 TSMC_233 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_25 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 
+ TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 
+ TSMC_1013 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_195 TSMC_196 
+ TSMC_1018 TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 
+ TSMC_1024 TSMC_1025 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 
+ TSMC_1031 TSMC_1032 TSMC_1033 TSMC_61 TSMC_93 TSMC_125 TSMC_157 
+ TSMC_213 TSMC_214 VDDI VSSI TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_26 TSMC_1034 TSMC_1035 TSMC_1036 TSMC_1037 TSMC_1038 
+ TSMC_1039 TSMC_1040 TSMC_1041 TSMC_1042 TSMC_1043 TSMC_1044 
+ TSMC_1045 TSMC_1046 TSMC_1047 TSMC_1048 TSMC_1049 TSMC_195 TSMC_196 
+ TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 TSMC_1062 
+ TSMC_1063 TSMC_1064 TSMC_1065 TSMC_62 TSMC_94 TSMC_126 TSMC_158 
+ TSMC_213 TSMC_214 VDDI VSSI TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_27 TSMC_1066 TSMC_1067 TSMC_1068 TSMC_1069 TSMC_1070 
+ TSMC_1071 TSMC_1072 TSMC_1073 TSMC_1074 TSMC_1075 TSMC_1076 
+ TSMC_1077 TSMC_1078 TSMC_1079 TSMC_1080 TSMC_1081 TSMC_195 TSMC_196 
+ TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 TSMC_1086 TSMC_1087 
+ TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 TSMC_1092 TSMC_1093 TSMC_1094 
+ TSMC_1095 TSMC_1096 TSMC_1097 TSMC_63 TSMC_95 TSMC_127 TSMC_159 
+ TSMC_213 TSMC_214 VDDI VSSI TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_28 TSMC_1098 TSMC_1099 TSMC_1100 TSMC_1101 TSMC_1102 
+ TSMC_1103 TSMC_1104 TSMC_1105 TSMC_1106 TSMC_1107 TSMC_1108 
+ TSMC_1109 TSMC_1110 TSMC_1111 TSMC_1112 TSMC_1113 TSMC_195 TSMC_196 
+ TSMC_1114 TSMC_1115 TSMC_1116 TSMC_1117 TSMC_1118 TSMC_1119 
+ TSMC_1120 TSMC_1121 TSMC_1122 TSMC_1123 TSMC_1124 TSMC_1125 TSMC_1126 
+ TSMC_1127 TSMC_1128 TSMC_1129 TSMC_64 TSMC_96 TSMC_128 TSMC_160 
+ TSMC_213 TSMC_214 VDDI VSSI TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_29 TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 
+ TSMC_1135 TSMC_1136 TSMC_1137 TSMC_1138 TSMC_1139 TSMC_1140 
+ TSMC_1141 TSMC_1142 TSMC_1143 TSMC_1144 TSMC_1145 TSMC_195 TSMC_196 
+ TSMC_1146 TSMC_1147 TSMC_1148 TSMC_1149 TSMC_1150 TSMC_1151 
+ TSMC_1152 TSMC_1153 TSMC_1154 TSMC_1155 TSMC_1156 TSMC_1157 TSMC_1158 
+ TSMC_1159 TSMC_1160 TSMC_1161 TSMC_65 TSMC_97 TSMC_129 TSMC_161 
+ TSMC_213 TSMC_214 VDDI VSSI TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_30 TSMC_1162 TSMC_1163 TSMC_1164 TSMC_1165 TSMC_1166 
+ TSMC_1167 TSMC_1168 TSMC_1169 TSMC_1170 TSMC_1171 TSMC_1172 
+ TSMC_1173 TSMC_1174 TSMC_1175 TSMC_1176 TSMC_1177 TSMC_195 TSMC_196 
+ TSMC_1178 TSMC_1179 TSMC_1180 TSMC_1181 TSMC_1182 TSMC_1183 
+ TSMC_1184 TSMC_1185 TSMC_1186 TSMC_1187 TSMC_1188 TSMC_1189 TSMC_1190 
+ TSMC_1191 TSMC_1192 TSMC_1193 TSMC_66 TSMC_98 TSMC_130 TSMC_162 
+ TSMC_213 TSMC_214 VDDI VSSI TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_31 TSMC_1194 TSMC_1195 TSMC_1196 TSMC_1197 TSMC_1198 
+ TSMC_1199 TSMC_1200 TSMC_1201 TSMC_1202 TSMC_1203 TSMC_1204 
+ TSMC_1205 TSMC_1206 TSMC_1207 TSMC_1208 TSMC_1209 TSMC_195 TSMC_196 
+ TSMC_1210 TSMC_1211 TSMC_1212 TSMC_1213 TSMC_1214 TSMC_1215 
+ TSMC_1216 TSMC_1217 TSMC_1218 TSMC_1219 TSMC_1220 TSMC_1221 TSMC_1222 
+ TSMC_1223 TSMC_1224 TSMC_1225 TSMC_67 TSMC_99 TSMC_131 TSMC_163 
+ TSMC_213 TSMC_214 VDDI VSSI TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 S1ALLSVTSW2000X20_LIO_M8_S 
XLCNT TSMC_195 TSMC_196 TSMC_1226 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 
+ TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 
+ TSMC_1227 TSMC_1228 TSMC_1229 TSMC_1230 TSMC_1231 TSMC_1232 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 
+ TSMC_233 TSMC_32 TSMC_33 TSMC_34 TSMC_1233 TSMC_1234 TSMC_35 
+ TSMC_1235 TSMC_1236 TSMC_1237 TSMC_1235 TSMC_165 TSMC_213 TSMC_214 
+ TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 TSMC_1238 VDDAI VDDHD 
+ VDDI TSMC_1239 TSMC_1235 VSSI TSMC_173 TSMC_215 TSMC_1240 TSMC_1241 
+ TSMC_1242 TSMC_1243 TSMC_1244 TSMC_1245 TSMC_1246 TSMC_1247 TSMC_174 
+ TSMC_1248 S1ALLSVTSW2000X20_LCTRL_M8_S 
XGTRK TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 TSMC_719 TSMC_720 
+ TSMC_721 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 TSMC_751 
+ TSMC_752 TSMC_753 TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_782 
+ TSMC_783 TSMC_784 TSMC_785 TSMC_810 TSMC_811 TSMC_812 TSMC_813 
+ TSMC_814 TSMC_815 TSMC_816 TSMC_817 TSMC_842 TSMC_843 TSMC_844 
+ TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_874 
+ TSMC_875 TSMC_876 TSMC_877 TSMC_878 TSMC_879 TSMC_880 TSMC_881 
+ TSMC_906 TSMC_907 TSMC_908 TSMC_909 TSMC_910 TSMC_911 TSMC_912 
+ TSMC_913 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 TSMC_943 
+ TSMC_944 TSMC_945 TSMC_970 TSMC_971 TSMC_972 TSMC_973 TSMC_974 
+ TSMC_975 TSMC_976 TSMC_977 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 
+ TSMC_1006 TSMC_1007 TSMC_1008 TSMC_1009 TSMC_1034 TSMC_1035 
+ TSMC_1036 TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 
+ TSMC_1066 TSMC_1067 TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 
+ TSMC_1072 TSMC_1073 TSMC_1098 TSMC_1099 TSMC_1100 TSMC_1101 
+ TSMC_1102 TSMC_1103 TSMC_1104 TSMC_1105 TSMC_1130 TSMC_1131 
+ TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 TSMC_1137 
+ TSMC_1162 TSMC_1163 TSMC_1164 TSMC_1165 TSMC_1166 TSMC_1167 
+ TSMC_1168 TSMC_1169 TSMC_1194 TSMC_1195 TSMC_1196 TSMC_1197 
+ TSMC_1198 TSMC_1199 TSMC_1200 TSMC_1201 TSMC_171 TSMC_1238 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 TSMC_1 
+ S1ALLSVTSW2000X20_GTRK_ARR 
XWLDV_256D TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_1505 TSMC_1506 TSMC_1227 
+ TSMC_1228 TSMC_1229 TSMC_1230 TSMC_1231 TSMC_1232 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_34 TSMC_164 
+ TSMC_165 TSMC_166 TSMC_168 TSMC_169 TSMC_1238 TSMC_1507 VDDHD VDDI VSSI 
+ TSMC_173 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 TSMC_1240 TSMC_1241 TSMC_1242 
+ TSMC_1243 TSMC_174 TSMC_1248 TSMC_175 TSMC_176 TSMC_177 TSMC_178 
+ S1ALLSVTSW2000X20_WLDV_F_DN 
XWLDV_256U TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_1505 TSMC_1506 TSMC_1227 
+ TSMC_1228 TSMC_1229 TSMC_1230 TSMC_1231 TSMC_1232 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_35 TSMC_164 
+ TSMC_165 TSMC_167 TSMC_168 TSMC_169 TSMC_1238 TSMC_1507 VDDHD VDDI VSSI 
+ TSMC_173 TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 
+ TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 
+ TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 
+ TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 
+ TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 
+ TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 
+ TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 
+ TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 
+ TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 
+ TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 TSMC_1244 TSMC_1245 
+ TSMC_1246 TSMC_1247 TSMC_174 TSMC_1248 TSMC_175 TSMC_176 TSMC_177 
+ TSMC_178 S1ALLSVTSW2000X20_WLDV_F 
XMCB_D0 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 
+ TSMC_204 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 
+ TSMC_185 TSMC_186 TSMC_36 TSMC_68 TSMC_100 TSMC_132 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 
+ TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 
+ TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 TSMC_1339 
+ TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1377 
+ TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 
+ TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 
+ TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U0 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 
+ TSMC_212 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_36 TSMC_68 TSMC_100 TSMC_132 VDDAI VDDI VSSI TSMC_1508 
+ TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 TSMC_1527 
+ TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 TSMC_1571 
+ TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 TSMC_1590 
+ TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 TSMC_1634 
+ TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 TSMC_1653 
+ TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 
+ TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 TSMC_1716 
+ TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 TSMC_1760 
+ TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D1 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 
+ TSMC_257 TSMC_234 TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 
+ TSMC_240 TSMC_241 TSMC_37 TSMC_69 TSMC_101 TSMC_133 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U1 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 
+ TSMC_265 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_37 TSMC_69 TSMC_101 TSMC_133 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D2 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 
+ TSMC_289 TSMC_266 TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 
+ TSMC_272 TSMC_273 TSMC_38 TSMC_70 TSMC_102 TSMC_134 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U2 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 
+ TSMC_297 TSMC_274 TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 
+ TSMC_280 TSMC_281 TSMC_38 TSMC_70 TSMC_102 TSMC_134 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D3 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 TSMC_319 TSMC_320 
+ TSMC_321 TSMC_298 TSMC_299 TSMC_300 TSMC_301 TSMC_302 TSMC_303 
+ TSMC_304 TSMC_305 TSMC_39 TSMC_71 TSMC_103 TSMC_135 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U3 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_326 TSMC_327 TSMC_328 
+ TSMC_329 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 
+ TSMC_312 TSMC_313 TSMC_39 TSMC_71 TSMC_103 TSMC_135 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D4 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 TSMC_351 TSMC_352 
+ TSMC_353 TSMC_330 TSMC_331 TSMC_332 TSMC_333 TSMC_334 TSMC_335 
+ TSMC_336 TSMC_337 TSMC_40 TSMC_72 TSMC_104 TSMC_136 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U4 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_358 TSMC_359 TSMC_360 
+ TSMC_361 TSMC_338 TSMC_339 TSMC_340 TSMC_341 TSMC_342 TSMC_343 
+ TSMC_344 TSMC_345 TSMC_40 TSMC_72 TSMC_104 TSMC_136 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D5 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 TSMC_383 TSMC_384 
+ TSMC_385 TSMC_362 TSMC_363 TSMC_364 TSMC_365 TSMC_366 TSMC_367 
+ TSMC_368 TSMC_369 TSMC_41 TSMC_73 TSMC_105 TSMC_137 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U5 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_390 TSMC_391 TSMC_392 
+ TSMC_393 TSMC_370 TSMC_371 TSMC_372 TSMC_373 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_41 TSMC_73 TSMC_105 TSMC_137 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D6 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 TSMC_415 TSMC_416 
+ TSMC_417 TSMC_394 TSMC_395 TSMC_396 TSMC_397 TSMC_398 TSMC_399 
+ TSMC_400 TSMC_401 TSMC_42 TSMC_74 TSMC_106 TSMC_138 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U6 TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_422 TSMC_423 TSMC_424 
+ TSMC_425 TSMC_402 TSMC_403 TSMC_404 TSMC_405 TSMC_406 TSMC_407 
+ TSMC_408 TSMC_409 TSMC_42 TSMC_74 TSMC_106 TSMC_138 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D7 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 TSMC_447 TSMC_448 
+ TSMC_449 TSMC_426 TSMC_427 TSMC_428 TSMC_429 TSMC_430 TSMC_431 
+ TSMC_432 TSMC_433 TSMC_43 TSMC_75 TSMC_107 TSMC_139 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U7 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_454 TSMC_455 TSMC_456 
+ TSMC_457 TSMC_434 TSMC_435 TSMC_436 TSMC_437 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_43 TSMC_75 TSMC_107 TSMC_139 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D8 TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 TSMC_479 TSMC_480 
+ TSMC_481 TSMC_458 TSMC_459 TSMC_460 TSMC_461 TSMC_462 TSMC_463 
+ TSMC_464 TSMC_465 TSMC_44 TSMC_76 TSMC_108 TSMC_140 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U8 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_486 TSMC_487 TSMC_488 
+ TSMC_489 TSMC_466 TSMC_467 TSMC_468 TSMC_469 TSMC_470 TSMC_471 
+ TSMC_472 TSMC_473 TSMC_44 TSMC_76 TSMC_108 TSMC_140 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D9 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 TSMC_511 TSMC_512 
+ TSMC_513 TSMC_490 TSMC_491 TSMC_492 TSMC_493 TSMC_494 TSMC_495 
+ TSMC_496 TSMC_497 TSMC_45 TSMC_77 TSMC_109 TSMC_141 VDDAI VDDI VSSI TSMC_1249 
+ TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 
+ TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 
+ TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 
+ TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 
+ TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 
+ TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 
+ TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 
+ TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U9 TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_518 TSMC_519 TSMC_520 
+ TSMC_521 TSMC_498 TSMC_499 TSMC_500 TSMC_501 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_45 TSMC_77 TSMC_109 TSMC_141 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D10 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 TSMC_543 
+ TSMC_544 TSMC_545 TSMC_522 TSMC_523 TSMC_524 TSMC_525 TSMC_526 
+ TSMC_527 TSMC_528 TSMC_529 TSMC_46 TSMC_78 TSMC_110 TSMC_142 VDDAI VDDI VSSI 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U10 TSMC_546 TSMC_547 TSMC_548 TSMC_549 TSMC_550 TSMC_551 
+ TSMC_552 TSMC_553 TSMC_530 TSMC_531 TSMC_532 TSMC_533 TSMC_534 
+ TSMC_535 TSMC_536 TSMC_537 TSMC_46 TSMC_78 TSMC_110 TSMC_142 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 
+ TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 
+ TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 
+ TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 
+ TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 
+ TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 
+ TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 
+ TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 
+ TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 
+ TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D11 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 TSMC_575 
+ TSMC_576 TSMC_577 TSMC_554 TSMC_555 TSMC_556 TSMC_557 TSMC_558 
+ TSMC_559 TSMC_560 TSMC_561 TSMC_47 TSMC_79 TSMC_111 TSMC_143 VDDAI VDDI VSSI 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U11 TSMC_578 TSMC_579 TSMC_580 TSMC_581 TSMC_582 TSMC_583 
+ TSMC_584 TSMC_585 TSMC_562 TSMC_563 TSMC_564 TSMC_565 TSMC_566 
+ TSMC_567 TSMC_568 TSMC_569 TSMC_47 TSMC_79 TSMC_111 TSMC_143 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 
+ TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 
+ TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 
+ TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 
+ TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 
+ TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 
+ TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 
+ TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 
+ TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 
+ TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D12 TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 TSMC_607 
+ TSMC_608 TSMC_609 TSMC_586 TSMC_587 TSMC_588 TSMC_589 TSMC_590 
+ TSMC_591 TSMC_592 TSMC_593 TSMC_48 TSMC_80 TSMC_112 TSMC_144 VDDAI VDDI 
+ VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 TSMC_1255 
+ TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 TSMC_1268 
+ TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 TSMC_1274 
+ TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 
+ TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 TSMC_1287 
+ TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 TSMC_1300 
+ TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 TSMC_1313 
+ TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 TSMC_1319 
+ TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 TSMC_1332 
+ TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 TSMC_1345 
+ TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 TSMC_1351 
+ TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 TSMC_1364 
+ TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 TSMC_1370 
+ TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 TSMC_1383 
+ TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 TSMC_1389 
+ TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 TSMC_1395 
+ TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 TSMC_1408 
+ TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 TSMC_1414 
+ TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 TSMC_1427 
+ TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 TSMC_1433 
+ TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 TSMC_1446 
+ TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 TSMC_1452 
+ TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 TSMC_1458 
+ TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 TSMC_1471 
+ TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 TSMC_1477 
+ TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 TSMC_1490 
+ TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 TSMC_1496 
+ TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U12 TSMC_610 TSMC_611 TSMC_612 TSMC_613 TSMC_614 TSMC_615 
+ TSMC_616 TSMC_617 TSMC_594 TSMC_595 TSMC_596 TSMC_597 TSMC_598 
+ TSMC_599 TSMC_600 TSMC_601 TSMC_48 TSMC_80 TSMC_112 TSMC_144 VDDAI VDDI 
+ VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 
+ TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 
+ TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D13 TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 TSMC_639 
+ TSMC_640 TSMC_641 TSMC_618 TSMC_619 TSMC_620 TSMC_621 TSMC_622 
+ TSMC_623 TSMC_624 TSMC_625 TSMC_49 TSMC_81 TSMC_113 TSMC_145 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U13 TSMC_642 TSMC_643 TSMC_644 TSMC_645 TSMC_646 TSMC_647 
+ TSMC_648 TSMC_649 TSMC_626 TSMC_627 TSMC_628 TSMC_629 TSMC_630 
+ TSMC_631 TSMC_632 TSMC_633 TSMC_49 TSMC_81 TSMC_113 TSMC_145 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D14 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 TSMC_671 
+ TSMC_672 TSMC_673 TSMC_650 TSMC_651 TSMC_652 TSMC_653 TSMC_654 
+ TSMC_655 TSMC_656 TSMC_657 TSMC_50 TSMC_82 TSMC_114 TSMC_146 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U14 TSMC_674 TSMC_675 TSMC_676 TSMC_677 TSMC_678 TSMC_679 
+ TSMC_680 TSMC_681 TSMC_658 TSMC_659 TSMC_660 TSMC_661 TSMC_662 
+ TSMC_663 TSMC_664 TSMC_665 TSMC_50 TSMC_82 TSMC_114 TSMC_146 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D15 TSMC_698 TSMC_699 TSMC_700 TSMC_701 TSMC_702 TSMC_703 
+ TSMC_704 TSMC_705 TSMC_682 TSMC_683 TSMC_684 TSMC_685 TSMC_686 
+ TSMC_687 TSMC_688 TSMC_689 TSMC_51 TSMC_83 TSMC_115 TSMC_147 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U15 TSMC_706 TSMC_707 TSMC_708 TSMC_709 TSMC_710 TSMC_711 
+ TSMC_712 TSMC_713 TSMC_690 TSMC_691 TSMC_692 TSMC_693 TSMC_694 
+ TSMC_695 TSMC_696 TSMC_697 TSMC_51 TSMC_83 TSMC_115 TSMC_147 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D16 TSMC_730 TSMC_731 TSMC_732 TSMC_733 TSMC_734 TSMC_735 
+ TSMC_736 TSMC_737 TSMC_714 TSMC_715 TSMC_716 TSMC_717 TSMC_718 
+ TSMC_719 TSMC_720 TSMC_721 TSMC_52 TSMC_84 TSMC_116 TSMC_148 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U16 TSMC_738 TSMC_739 TSMC_740 TSMC_741 TSMC_742 TSMC_743 
+ TSMC_744 TSMC_745 TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_726 
+ TSMC_727 TSMC_728 TSMC_729 TSMC_52 TSMC_84 TSMC_116 TSMC_148 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D17 TSMC_762 TSMC_763 TSMC_764 TSMC_765 TSMC_766 TSMC_767 
+ TSMC_768 TSMC_769 TSMC_746 TSMC_747 TSMC_748 TSMC_749 TSMC_750 
+ TSMC_751 TSMC_752 TSMC_753 TSMC_53 TSMC_85 TSMC_117 TSMC_149 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U17 TSMC_770 TSMC_771 TSMC_772 TSMC_773 TSMC_774 TSMC_775 
+ TSMC_776 TSMC_777 TSMC_754 TSMC_755 TSMC_756 TSMC_757 TSMC_758 
+ TSMC_759 TSMC_760 TSMC_761 TSMC_53 TSMC_85 TSMC_117 TSMC_149 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D18 TSMC_794 TSMC_795 TSMC_796 TSMC_797 TSMC_798 TSMC_799 
+ TSMC_800 TSMC_801 TSMC_778 TSMC_779 TSMC_780 TSMC_781 TSMC_782 
+ TSMC_783 TSMC_784 TSMC_785 TSMC_54 TSMC_86 TSMC_118 TSMC_150 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U18 TSMC_802 TSMC_803 TSMC_804 TSMC_805 TSMC_806 TSMC_807 
+ TSMC_808 TSMC_809 TSMC_786 TSMC_787 TSMC_788 TSMC_789 TSMC_790 
+ TSMC_791 TSMC_792 TSMC_793 TSMC_54 TSMC_86 TSMC_118 TSMC_150 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D19 TSMC_826 TSMC_827 TSMC_828 TSMC_829 TSMC_830 TSMC_831 
+ TSMC_832 TSMC_833 TSMC_810 TSMC_811 TSMC_812 TSMC_813 TSMC_814 
+ TSMC_815 TSMC_816 TSMC_817 TSMC_55 TSMC_87 TSMC_119 TSMC_151 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U19 TSMC_834 TSMC_835 TSMC_836 TSMC_837 TSMC_838 TSMC_839 
+ TSMC_840 TSMC_841 TSMC_818 TSMC_819 TSMC_820 TSMC_821 TSMC_822 
+ TSMC_823 TSMC_824 TSMC_825 TSMC_55 TSMC_87 TSMC_119 TSMC_151 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D20 TSMC_858 TSMC_859 TSMC_860 TSMC_861 TSMC_862 TSMC_863 
+ TSMC_864 TSMC_865 TSMC_842 TSMC_843 TSMC_844 TSMC_845 TSMC_846 
+ TSMC_847 TSMC_848 TSMC_849 TSMC_56 TSMC_88 TSMC_120 TSMC_152 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U20 TSMC_866 TSMC_867 TSMC_868 TSMC_869 TSMC_870 TSMC_871 
+ TSMC_872 TSMC_873 TSMC_850 TSMC_851 TSMC_852 TSMC_853 TSMC_854 
+ TSMC_855 TSMC_856 TSMC_857 TSMC_56 TSMC_88 TSMC_120 TSMC_152 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D21 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 TSMC_895 
+ TSMC_896 TSMC_897 TSMC_874 TSMC_875 TSMC_876 TSMC_877 TSMC_878 
+ TSMC_879 TSMC_880 TSMC_881 TSMC_57 TSMC_89 TSMC_121 TSMC_153 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U21 TSMC_898 TSMC_899 TSMC_900 TSMC_901 TSMC_902 TSMC_903 
+ TSMC_904 TSMC_905 TSMC_882 TSMC_883 TSMC_884 TSMC_885 TSMC_886 
+ TSMC_887 TSMC_888 TSMC_889 TSMC_57 TSMC_89 TSMC_121 TSMC_153 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D22 TSMC_922 TSMC_923 TSMC_924 TSMC_925 TSMC_926 TSMC_927 
+ TSMC_928 TSMC_929 TSMC_906 TSMC_907 TSMC_908 TSMC_909 TSMC_910 
+ TSMC_911 TSMC_912 TSMC_913 TSMC_58 TSMC_90 TSMC_122 TSMC_154 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U22 TSMC_930 TSMC_931 TSMC_932 TSMC_933 TSMC_934 TSMC_935 
+ TSMC_936 TSMC_937 TSMC_914 TSMC_915 TSMC_916 TSMC_917 TSMC_918 
+ TSMC_919 TSMC_920 TSMC_921 TSMC_58 TSMC_90 TSMC_122 TSMC_154 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D23 TSMC_954 TSMC_955 TSMC_956 TSMC_957 TSMC_958 TSMC_959 
+ TSMC_960 TSMC_961 TSMC_938 TSMC_939 TSMC_940 TSMC_941 TSMC_942 
+ TSMC_943 TSMC_944 TSMC_945 TSMC_59 TSMC_91 TSMC_123 TSMC_155 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U23 TSMC_962 TSMC_963 TSMC_964 TSMC_965 TSMC_966 TSMC_967 
+ TSMC_968 TSMC_969 TSMC_946 TSMC_947 TSMC_948 TSMC_949 TSMC_950 
+ TSMC_951 TSMC_952 TSMC_953 TSMC_59 TSMC_91 TSMC_123 TSMC_155 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D24 TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 TSMC_991 
+ TSMC_992 TSMC_993 TSMC_970 TSMC_971 TSMC_972 TSMC_973 TSMC_974 
+ TSMC_975 TSMC_976 TSMC_977 TSMC_60 TSMC_92 TSMC_124 TSMC_156 VDDAI 
+ VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 TSMC_1504 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U24 TSMC_994 TSMC_995 TSMC_996 TSMC_997 TSMC_998 TSMC_999 
+ TSMC_1000 TSMC_1001 TSMC_978 TSMC_979 TSMC_980 TSMC_981 TSMC_982 
+ TSMC_983 TSMC_984 TSMC_985 TSMC_60 TSMC_92 TSMC_124 TSMC_156 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D25 TSMC_1018 TSMC_1019 TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 
+ TSMC_1024 TSMC_1025 TSMC_1002 TSMC_1003 TSMC_1004 TSMC_1005 
+ TSMC_1006 TSMC_1007 TSMC_1008 TSMC_1009 TSMC_61 TSMC_93 TSMC_125 
+ TSMC_157 VDDAI VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U25 TSMC_1026 TSMC_1027 TSMC_1028 TSMC_1029 TSMC_1030 TSMC_1031 
+ TSMC_1032 TSMC_1033 TSMC_1010 TSMC_1011 TSMC_1012 TSMC_1013 
+ TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_61 TSMC_93 TSMC_125 
+ TSMC_157 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D26 TSMC_1050 TSMC_1051 TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 
+ TSMC_1056 TSMC_1057 TSMC_1034 TSMC_1035 TSMC_1036 TSMC_1037 
+ TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 TSMC_62 TSMC_94 TSMC_126 
+ TSMC_158 VDDAI VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U26 TSMC_1058 TSMC_1059 TSMC_1060 TSMC_1061 TSMC_1062 TSMC_1063 
+ TSMC_1064 TSMC_1065 TSMC_1042 TSMC_1043 TSMC_1044 TSMC_1045 
+ TSMC_1046 TSMC_1047 TSMC_1048 TSMC_1049 TSMC_62 TSMC_94 TSMC_126 
+ TSMC_158 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D27 TSMC_1082 TSMC_1083 TSMC_1084 TSMC_1085 TSMC_1086 TSMC_1087 
+ TSMC_1088 TSMC_1089 TSMC_1066 TSMC_1067 TSMC_1068 TSMC_1069 
+ TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 TSMC_63 TSMC_95 TSMC_127 
+ TSMC_159 VDDAI VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U27 TSMC_1090 TSMC_1091 TSMC_1092 TSMC_1093 TSMC_1094 TSMC_1095 
+ TSMC_1096 TSMC_1097 TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 
+ TSMC_1078 TSMC_1079 TSMC_1080 TSMC_1081 TSMC_63 TSMC_95 TSMC_127 
+ TSMC_159 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D28 TSMC_1114 TSMC_1115 TSMC_1116 TSMC_1117 TSMC_1118 TSMC_1119 
+ TSMC_1120 TSMC_1121 TSMC_1098 TSMC_1099 TSMC_1100 TSMC_1101 
+ TSMC_1102 TSMC_1103 TSMC_1104 TSMC_1105 TSMC_64 TSMC_96 TSMC_128 
+ TSMC_160 VDDAI VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U28 TSMC_1122 TSMC_1123 TSMC_1124 TSMC_1125 TSMC_1126 TSMC_1127 
+ TSMC_1128 TSMC_1129 TSMC_1106 TSMC_1107 TSMC_1108 TSMC_1109 
+ TSMC_1110 TSMC_1111 TSMC_1112 TSMC_1113 TSMC_64 TSMC_96 TSMC_128 
+ TSMC_160 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D29 TSMC_1146 TSMC_1147 TSMC_1148 TSMC_1149 TSMC_1150 TSMC_1151 
+ TSMC_1152 TSMC_1153 TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 
+ TSMC_1134 TSMC_1135 TSMC_1136 TSMC_1137 TSMC_65 TSMC_97 TSMC_129 
+ TSMC_161 VDDAI VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U29 TSMC_1154 TSMC_1155 TSMC_1156 TSMC_1157 TSMC_1158 TSMC_1159 
+ TSMC_1160 TSMC_1161 TSMC_1138 TSMC_1139 TSMC_1140 TSMC_1141 
+ TSMC_1142 TSMC_1143 TSMC_1144 TSMC_1145 TSMC_65 TSMC_97 TSMC_129 
+ TSMC_161 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D30 TSMC_1178 TSMC_1179 TSMC_1180 TSMC_1181 TSMC_1182 TSMC_1183 
+ TSMC_1184 TSMC_1185 TSMC_1162 TSMC_1163 TSMC_1164 TSMC_1165 
+ TSMC_1166 TSMC_1167 TSMC_1168 TSMC_1169 TSMC_66 TSMC_98 TSMC_130 
+ TSMC_162 VDDAI VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U30 TSMC_1186 TSMC_1187 TSMC_1188 TSMC_1189 TSMC_1190 TSMC_1191 
+ TSMC_1192 TSMC_1193 TSMC_1170 TSMC_1171 TSMC_1172 TSMC_1173 
+ TSMC_1174 TSMC_1175 TSMC_1176 TSMC_1177 TSMC_66 TSMC_98 TSMC_130 
+ TSMC_162 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D31 TSMC_1210 TSMC_1211 TSMC_1212 TSMC_1213 TSMC_1214 TSMC_1215 
+ TSMC_1216 TSMC_1217 TSMC_1194 TSMC_1195 TSMC_1196 TSMC_1197 
+ TSMC_1198 TSMC_1199 TSMC_1200 TSMC_1201 TSMC_67 TSMC_99 TSMC_131 
+ TSMC_163 VDDAI VDDI VSSI TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1504 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U31 TSMC_1218 TSMC_1219 TSMC_1220 TSMC_1221 TSMC_1222 TSMC_1223 
+ TSMC_1224 TSMC_1225 TSMC_1202 TSMC_1203 TSMC_1204 TSMC_1205 
+ TSMC_1206 TSMC_1207 TSMC_1208 TSMC_1209 TSMC_67 TSMC_99 TSMC_131 
+ TSMC_163 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
.ENDS

.SUBCKT S1ALLSVTSW2000X20_BANK_F TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 VDDAI VDDHD VDDI VSSI TSMC_171 TSMC_172 TSMC_173 TSMC_174 
XLIO_M8_S_AL_0 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 
+ TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 
+ TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 
+ TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 
+ TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_35 
+ TSMC_67 TSMC_99 TSMC_131 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_1 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_191 TSMC_192 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 
+ TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 TSMC_36 
+ TSMC_68 TSMC_100 TSMC_132 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_2 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 
+ TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 
+ TSMC_275 TSMC_276 TSMC_277 TSMC_191 TSMC_192 TSMC_278 TSMC_279 
+ TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 TSMC_285 TSMC_286 
+ TSMC_287 TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 TSMC_37 
+ TSMC_69 TSMC_101 TSMC_133 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_3 TSMC_294 TSMC_295 TSMC_296 TSMC_297 TSMC_298 TSMC_299 
+ TSMC_300 TSMC_301 TSMC_302 TSMC_303 TSMC_304 TSMC_305 TSMC_306 
+ TSMC_307 TSMC_308 TSMC_309 TSMC_191 TSMC_192 TSMC_310 TSMC_311 
+ TSMC_312 TSMC_313 TSMC_314 TSMC_315 TSMC_316 TSMC_317 TSMC_318 
+ TSMC_319 TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 TSMC_325 TSMC_38 
+ TSMC_70 TSMC_102 TSMC_134 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_4 TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 
+ TSMC_332 TSMC_333 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 
+ TSMC_339 TSMC_340 TSMC_341 TSMC_191 TSMC_192 TSMC_342 TSMC_343 
+ TSMC_344 TSMC_345 TSMC_346 TSMC_347 TSMC_348 TSMC_349 TSMC_350 
+ TSMC_351 TSMC_352 TSMC_353 TSMC_354 TSMC_355 TSMC_356 TSMC_357 TSMC_39 
+ TSMC_71 TSMC_103 TSMC_135 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_5 TSMC_358 TSMC_359 TSMC_360 TSMC_361 TSMC_362 TSMC_363 
+ TSMC_364 TSMC_365 TSMC_366 TSMC_367 TSMC_368 TSMC_369 TSMC_370 
+ TSMC_371 TSMC_372 TSMC_373 TSMC_191 TSMC_192 TSMC_374 TSMC_375 
+ TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 TSMC_381 TSMC_382 
+ TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 TSMC_389 TSMC_40 
+ TSMC_72 TSMC_104 TSMC_136 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_6 TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 
+ TSMC_396 TSMC_397 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 
+ TSMC_403 TSMC_404 TSMC_405 TSMC_191 TSMC_192 TSMC_406 TSMC_407 
+ TSMC_408 TSMC_409 TSMC_410 TSMC_411 TSMC_412 TSMC_413 TSMC_414 
+ TSMC_415 TSMC_416 TSMC_417 TSMC_418 TSMC_419 TSMC_420 TSMC_421 TSMC_41 
+ TSMC_73 TSMC_105 TSMC_137 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_7 TSMC_422 TSMC_423 TSMC_424 TSMC_425 TSMC_426 TSMC_427 
+ TSMC_428 TSMC_429 TSMC_430 TSMC_431 TSMC_432 TSMC_433 TSMC_434 
+ TSMC_435 TSMC_436 TSMC_437 TSMC_191 TSMC_192 TSMC_438 TSMC_439 
+ TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 TSMC_445 TSMC_446 
+ TSMC_447 TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 TSMC_453 TSMC_42 
+ TSMC_74 TSMC_106 TSMC_138 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_8 TSMC_454 TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 
+ TSMC_460 TSMC_461 TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 
+ TSMC_467 TSMC_468 TSMC_469 TSMC_191 TSMC_192 TSMC_470 TSMC_471 
+ TSMC_472 TSMC_473 TSMC_474 TSMC_475 TSMC_476 TSMC_477 TSMC_478 
+ TSMC_479 TSMC_480 TSMC_481 TSMC_482 TSMC_483 TSMC_484 TSMC_485 TSMC_43 
+ TSMC_75 TSMC_107 TSMC_139 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_9 TSMC_486 TSMC_487 TSMC_488 TSMC_489 TSMC_490 TSMC_491 
+ TSMC_492 TSMC_493 TSMC_494 TSMC_495 TSMC_496 TSMC_497 TSMC_498 
+ TSMC_499 TSMC_500 TSMC_501 TSMC_191 TSMC_192 TSMC_502 TSMC_503 
+ TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 TSMC_509 TSMC_510 
+ TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 TSMC_517 TSMC_44 
+ TSMC_76 TSMC_108 TSMC_140 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_AL_10 TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 TSMC_523 
+ TSMC_524 TSMC_525 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 
+ TSMC_531 TSMC_532 TSMC_533 TSMC_191 TSMC_192 TSMC_534 TSMC_535 
+ TSMC_536 TSMC_537 TSMC_538 TSMC_539 TSMC_540 TSMC_541 TSMC_542 
+ TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 TSMC_548 TSMC_549 
+ TSMC_45 TSMC_77 TSMC_109 TSMC_141 TSMC_209 TSMC_210 VDDI VSSI 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_ABL_11 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 TSMC_555 
+ TSMC_556 TSMC_557 TSMC_558 TSMC_559 TSMC_560 TSMC_561 TSMC_562 
+ TSMC_563 TSMC_564 TSMC_565 TSMC_191 TSMC_192 TSMC_566 TSMC_567 
+ TSMC_568 TSMC_569 TSMC_570 TSMC_571 TSMC_572 TSMC_573 TSMC_574 
+ TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 TSMC_580 TSMC_581 
+ TSMC_46 TSMC_78 TSMC_110 TSMC_142 TSMC_209 TSMC_210 VDDI VSSI 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CL_12 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 TSMC_587 
+ TSMC_588 TSMC_589 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_191 TSMC_192 TSMC_598 TSMC_599 
+ TSMC_600 TSMC_601 TSMC_602 TSMC_603 TSMC_604 TSMC_605 TSMC_606 
+ TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 TSMC_612 TSMC_613 
+ TSMC_47 TSMC_79 TSMC_111 TSMC_143 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CL_13 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 TSMC_619 
+ TSMC_620 TSMC_621 TSMC_622 TSMC_623 TSMC_624 TSMC_625 TSMC_626 
+ TSMC_627 TSMC_628 TSMC_629 TSMC_191 TSMC_192 TSMC_630 TSMC_631 
+ TSMC_632 TSMC_633 TSMC_634 TSMC_635 TSMC_636 TSMC_637 TSMC_638 
+ TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 TSMC_644 TSMC_645 
+ TSMC_48 TSMC_80 TSMC_112 TSMC_144 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CL_14 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 TSMC_651 
+ TSMC_652 TSMC_653 TSMC_654 TSMC_655 TSMC_656 TSMC_657 TSMC_658 
+ TSMC_659 TSMC_660 TSMC_661 TSMC_191 TSMC_192 TSMC_662 TSMC_663 
+ TSMC_664 TSMC_665 TSMC_666 TSMC_667 TSMC_668 TSMC_669 TSMC_670 
+ TSMC_671 TSMC_672 TSMC_673 TSMC_674 TSMC_675 TSMC_676 TSMC_677 
+ TSMC_49 TSMC_81 TSMC_113 TSMC_145 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CBL_L_15 TSMC_678 TSMC_679 TSMC_680 TSMC_681 TSMC_682 
+ TSMC_683 TSMC_684 TSMC_685 TSMC_686 TSMC_687 TSMC_688 TSMC_689 
+ TSMC_690 TSMC_691 TSMC_692 TSMC_693 TSMC_191 TSMC_192 TSMC_694 
+ TSMC_695 TSMC_696 TSMC_697 TSMC_698 TSMC_699 TSMC_700 TSMC_701 
+ TSMC_702 TSMC_703 TSMC_704 TSMC_705 TSMC_706 TSMC_707 TSMC_708 
+ TSMC_709 TSMC_50 TSMC_82 TSMC_114 TSMC_146 TSMC_209 TSMC_210 VDDI VSSI 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_CBL_R_16 TSMC_710 TSMC_711 TSMC_712 TSMC_713 TSMC_714 
+ TSMC_715 TSMC_716 TSMC_717 TSMC_718 TSMC_719 TSMC_720 TSMC_721 
+ TSMC_722 TSMC_723 TSMC_724 TSMC_725 TSMC_191 TSMC_192 TSMC_726 
+ TSMC_727 TSMC_728 TSMC_729 TSMC_730 TSMC_731 TSMC_732 TSMC_733 
+ TSMC_734 TSMC_735 TSMC_736 TSMC_737 TSMC_738 TSMC_739 TSMC_740 
+ TSMC_741 TSMC_51 TSMC_83 TSMC_115 TSMC_147 TSMC_209 TSMC_210 VDDI VSSI 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_C_R_17 TSMC_742 TSMC_743 TSMC_744 TSMC_745 TSMC_746 TSMC_747 
+ TSMC_748 TSMC_749 TSMC_750 TSMC_751 TSMC_752 TSMC_753 TSMC_754 
+ TSMC_755 TSMC_756 TSMC_757 TSMC_191 TSMC_192 TSMC_758 TSMC_759 
+ TSMC_760 TSMC_761 TSMC_762 TSMC_763 TSMC_764 TSMC_765 TSMC_766 
+ TSMC_767 TSMC_768 TSMC_769 TSMC_770 TSMC_771 TSMC_772 TSMC_773 
+ TSMC_52 TSMC_84 TSMC_116 TSMC_148 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_C_R_18 TSMC_774 TSMC_775 TSMC_776 TSMC_777 TSMC_778 TSMC_779 
+ TSMC_780 TSMC_781 TSMC_782 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ TSMC_787 TSMC_788 TSMC_789 TSMC_191 TSMC_192 TSMC_790 TSMC_791 
+ TSMC_792 TSMC_793 TSMC_794 TSMC_795 TSMC_796 TSMC_797 TSMC_798 
+ TSMC_799 TSMC_800 TSMC_801 TSMC_802 TSMC_803 TSMC_804 TSMC_805 
+ TSMC_53 TSMC_85 TSMC_117 TSMC_149 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_C_R_19 TSMC_806 TSMC_807 TSMC_808 TSMC_809 TSMC_810 TSMC_811 
+ TSMC_812 TSMC_813 TSMC_814 TSMC_815 TSMC_816 TSMC_817 TSMC_818 
+ TSMC_819 TSMC_820 TSMC_821 TSMC_191 TSMC_192 TSMC_822 TSMC_823 
+ TSMC_824 TSMC_825 TSMC_826 TSMC_827 TSMC_828 TSMC_829 TSMC_830 
+ TSMC_831 TSMC_832 TSMC_833 TSMC_834 TSMC_835 TSMC_836 TSMC_837 
+ TSMC_54 TSMC_86 TSMC_118 TSMC_150 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_ABL_R_20 TSMC_838 TSMC_839 TSMC_840 TSMC_841 TSMC_842 
+ TSMC_843 TSMC_844 TSMC_845 TSMC_846 TSMC_847 TSMC_848 TSMC_849 
+ TSMC_850 TSMC_851 TSMC_852 TSMC_853 TSMC_191 TSMC_192 TSMC_854 
+ TSMC_855 TSMC_856 TSMC_857 TSMC_858 TSMC_859 TSMC_860 TSMC_861 
+ TSMC_862 TSMC_863 TSMC_864 TSMC_865 TSMC_866 TSMC_867 TSMC_868 
+ TSMC_869 TSMC_55 TSMC_87 TSMC_119 TSMC_151 TSMC_209 TSMC_210 VDDI VSSI 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 
+ TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 
+ TSMC_225 TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_21 TSMC_870 TSMC_871 TSMC_872 TSMC_873 TSMC_874 TSMC_875 
+ TSMC_876 TSMC_877 TSMC_878 TSMC_879 TSMC_880 TSMC_881 TSMC_882 
+ TSMC_883 TSMC_884 TSMC_885 TSMC_191 TSMC_192 TSMC_886 TSMC_887 
+ TSMC_888 TSMC_889 TSMC_890 TSMC_891 TSMC_892 TSMC_893 TSMC_894 
+ TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 TSMC_900 TSMC_901 
+ TSMC_56 TSMC_88 TSMC_120 TSMC_152 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_22 TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 TSMC_907 
+ TSMC_908 TSMC_909 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 
+ TSMC_915 TSMC_916 TSMC_917 TSMC_191 TSMC_192 TSMC_918 TSMC_919 
+ TSMC_920 TSMC_921 TSMC_922 TSMC_923 TSMC_924 TSMC_925 TSMC_926 
+ TSMC_927 TSMC_928 TSMC_929 TSMC_930 TSMC_931 TSMC_932 TSMC_933 
+ TSMC_57 TSMC_89 TSMC_121 TSMC_153 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_23 TSMC_934 TSMC_935 TSMC_936 TSMC_937 TSMC_938 TSMC_939 
+ TSMC_940 TSMC_941 TSMC_942 TSMC_943 TSMC_944 TSMC_945 TSMC_946 
+ TSMC_947 TSMC_948 TSMC_949 TSMC_191 TSMC_192 TSMC_950 TSMC_951 
+ TSMC_952 TSMC_953 TSMC_954 TSMC_955 TSMC_956 TSMC_957 TSMC_958 
+ TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 TSMC_964 TSMC_965 
+ TSMC_58 TSMC_90 TSMC_122 TSMC_154 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_24 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 TSMC_971 
+ TSMC_972 TSMC_973 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_191 TSMC_192 TSMC_982 TSMC_983 
+ TSMC_984 TSMC_985 TSMC_986 TSMC_987 TSMC_988 TSMC_989 TSMC_990 
+ TSMC_991 TSMC_992 TSMC_993 TSMC_994 TSMC_995 TSMC_996 TSMC_997 
+ TSMC_59 TSMC_91 TSMC_123 TSMC_155 TSMC_209 TSMC_210 VDDI VSSI TSMC_211 
+ TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 
+ TSMC_226 TSMC_227 TSMC_228 TSMC_229 
+ S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_25 TSMC_998 TSMC_999 TSMC_1000 TSMC_1001 TSMC_1002 
+ TSMC_1003 TSMC_1004 TSMC_1005 TSMC_1006 TSMC_1007 TSMC_1008 
+ TSMC_1009 TSMC_1010 TSMC_1011 TSMC_1012 TSMC_1013 TSMC_191 TSMC_192 
+ TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 TSMC_1019 
+ TSMC_1020 TSMC_1021 TSMC_1022 TSMC_1023 TSMC_1024 TSMC_1025 TSMC_1026 
+ TSMC_1027 TSMC_1028 TSMC_1029 TSMC_60 TSMC_92 TSMC_124 TSMC_156 
+ TSMC_209 TSMC_210 VDDI VSSI TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_26 TSMC_1030 TSMC_1031 TSMC_1032 TSMC_1033 TSMC_1034 
+ TSMC_1035 TSMC_1036 TSMC_1037 TSMC_1038 TSMC_1039 TSMC_1040 
+ TSMC_1041 TSMC_1042 TSMC_1043 TSMC_1044 TSMC_1045 TSMC_191 TSMC_192 
+ TSMC_1046 TSMC_1047 TSMC_1048 TSMC_1049 TSMC_1050 TSMC_1051 
+ TSMC_1052 TSMC_1053 TSMC_1054 TSMC_1055 TSMC_1056 TSMC_1057 TSMC_1058 
+ TSMC_1059 TSMC_1060 TSMC_1061 TSMC_61 TSMC_93 TSMC_125 TSMC_157 
+ TSMC_209 TSMC_210 VDDI VSSI TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_27 TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 TSMC_1066 
+ TSMC_1067 TSMC_1068 TSMC_1069 TSMC_1070 TSMC_1071 TSMC_1072 
+ TSMC_1073 TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_191 TSMC_192 
+ TSMC_1078 TSMC_1079 TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 
+ TSMC_1084 TSMC_1085 TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 
+ TSMC_1091 TSMC_1092 TSMC_1093 TSMC_62 TSMC_94 TSMC_126 TSMC_158 
+ TSMC_209 TSMC_210 VDDI VSSI TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_28 TSMC_1094 TSMC_1095 TSMC_1096 TSMC_1097 TSMC_1098 
+ TSMC_1099 TSMC_1100 TSMC_1101 TSMC_1102 TSMC_1103 TSMC_1104 
+ TSMC_1105 TSMC_1106 TSMC_1107 TSMC_1108 TSMC_1109 TSMC_191 TSMC_192 
+ TSMC_1110 TSMC_1111 TSMC_1112 TSMC_1113 TSMC_1114 TSMC_1115 
+ TSMC_1116 TSMC_1117 TSMC_1118 TSMC_1119 TSMC_1120 TSMC_1121 TSMC_1122 
+ TSMC_1123 TSMC_1124 TSMC_1125 TSMC_63 TSMC_95 TSMC_127 TSMC_159 
+ TSMC_209 TSMC_210 VDDI VSSI TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_29 TSMC_1126 TSMC_1127 TSMC_1128 TSMC_1129 TSMC_1130 
+ TSMC_1131 TSMC_1132 TSMC_1133 TSMC_1134 TSMC_1135 TSMC_1136 
+ TSMC_1137 TSMC_1138 TSMC_1139 TSMC_1140 TSMC_1141 TSMC_191 TSMC_192 
+ TSMC_1142 TSMC_1143 TSMC_1144 TSMC_1145 TSMC_1146 TSMC_1147 
+ TSMC_1148 TSMC_1149 TSMC_1150 TSMC_1151 TSMC_1152 TSMC_1153 TSMC_1154 
+ TSMC_1155 TSMC_1156 TSMC_1157 TSMC_64 TSMC_96 TSMC_128 TSMC_160 
+ TSMC_209 TSMC_210 VDDI VSSI TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_30 TSMC_1158 TSMC_1159 TSMC_1160 TSMC_1161 TSMC_1162 
+ TSMC_1163 TSMC_1164 TSMC_1165 TSMC_1166 TSMC_1167 TSMC_1168 
+ TSMC_1169 TSMC_1170 TSMC_1171 TSMC_1172 TSMC_1173 TSMC_191 TSMC_192 
+ TSMC_1174 TSMC_1175 TSMC_1176 TSMC_1177 TSMC_1178 TSMC_1179 
+ TSMC_1180 TSMC_1181 TSMC_1182 TSMC_1183 TSMC_1184 TSMC_1185 TSMC_1186 
+ TSMC_1187 TSMC_1188 TSMC_1189 TSMC_65 TSMC_97 TSMC_129 TSMC_161 
+ TSMC_209 TSMC_210 VDDI VSSI TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 S1ALLSVTSW2000X20_LIO_M8_S 
XLIO_M8_S_A_R_31 TSMC_1190 TSMC_1191 TSMC_1192 TSMC_1193 TSMC_1194 
+ TSMC_1195 TSMC_1196 TSMC_1197 TSMC_1198 TSMC_1199 TSMC_1200 
+ TSMC_1201 TSMC_1202 TSMC_1203 TSMC_1204 TSMC_1205 TSMC_191 TSMC_192 
+ TSMC_1206 TSMC_1207 TSMC_1208 TSMC_1209 TSMC_1210 TSMC_1211 
+ TSMC_1212 TSMC_1213 TSMC_1214 TSMC_1215 TSMC_1216 TSMC_1217 TSMC_1218 
+ TSMC_1219 TSMC_1220 TSMC_1221 TSMC_66 TSMC_98 TSMC_130 TSMC_162 
+ TSMC_209 TSMC_210 VDDI VSSI TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 
+ TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 TSMC_222 
+ TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 S1ALLSVTSW2000X20_LIO_M8_S 
XLCNT TSMC_191 TSMC_192 TSMC_1222 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 
+ TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 
+ TSMC_15 TSMC_16 TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 
+ TSMC_1223 TSMC_1224 TSMC_1225 TSMC_1226 TSMC_1227 TSMC_1228 TSMC_23 
+ TSMC_24 TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_214 
+ TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 TSMC_220 TSMC_221 
+ TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 TSMC_227 TSMC_228 
+ TSMC_229 TSMC_31 TSMC_32 TSMC_33 TSMC_1229 TSMC_1230 TSMC_34 
+ TSMC_1231 TSMC_1232 TSMC_1233 TSMC_1231 TSMC_164 TSMC_209 TSMC_210 
+ TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_1234 VDDAI VDDHD 
+ VDDI TSMC_1235 TSMC_1231 VSSI TSMC_171 TSMC_211 TSMC_1236 TSMC_1237 
+ TSMC_1238 TSMC_1239 TSMC_1240 TSMC_1241 TSMC_1242 TSMC_1243 TSMC_172 
+ TSMC_1244 S1ALLSVTSW2000X20_LCTRL_M8_S 
XWLDV_256D TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_1245 TSMC_1246 TSMC_1223 
+ TSMC_1224 TSMC_1225 TSMC_1226 TSMC_1227 TSMC_1228 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_33 TSMC_163 
+ TSMC_164 TSMC_165 TSMC_167 TSMC_168 TSMC_1234 TSMC_1247 VDDHD VDDI VSSI 
+ TSMC_171 TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 
+ TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 
+ TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 
+ TSMC_1272 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 
+ TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 
+ TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 
+ TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 
+ TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 
+ TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 
+ TSMC_1368 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 
+ TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 
+ TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 
+ TSMC_1412 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 
+ TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 
+ TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 
+ TSMC_1488 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 TSMC_1236 TSMC_1237 TSMC_1238 
+ TSMC_1239 TSMC_172 TSMC_1244 TSMC_173 TSMC_174 TSMC_1504 TSMC_1505 
+ S1ALLSVTSW2000X20_WLDV_F_DN 
XWLDV_256U TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_1245 TSMC_1246 TSMC_1223 
+ TSMC_1224 TSMC_1225 TSMC_1226 TSMC_1227 TSMC_1228 TSMC_23 TSMC_24 
+ TSMC_25 TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_1506 TSMC_163 
+ TSMC_164 TSMC_1507 TSMC_167 TSMC_168 TSMC_1234 TSMC_1247 VDDHD VDDI 
+ VSSI TSMC_171 TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 
+ TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 
+ TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 
+ TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 
+ TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 TSMC_1240 
+ TSMC_1241 TSMC_1242 TSMC_1243 TSMC_172 TSMC_1244 TSMC_173 TSMC_174 TSMC_1504 
+ TSMC_1505 S1ALLSVTSW2000X20_WLDV_F 
XMCB_D0 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 
+ TSMC_200 TSMC_175 TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 
+ TSMC_181 TSMC_182 TSMC_35 TSMC_67 TSMC_99 TSMC_131 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 TSMC_1261 
+ TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 TSMC_1306 
+ TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 TSMC_1338 
+ TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 TSMC_1376 
+ TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 TSMC_1439 
+ TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 TSMC_1502 
+ TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U0 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_183 TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 
+ TSMC_189 TSMC_190 TSMC_35 TSMC_67 TSMC_99 TSMC_131 VDDAI VDDI VSSI TSMC_1508 
+ TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 TSMC_1527 
+ TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 TSMC_1571 
+ TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 TSMC_1590 
+ TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 TSMC_1634 
+ TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 TSMC_1653 
+ TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 TSMC_1697 
+ TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 TSMC_1716 
+ TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 TSMC_1760 
+ TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D1 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 
+ TSMC_253 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 TSMC_235 
+ TSMC_236 TSMC_237 TSMC_36 TSMC_68 TSMC_100 TSMC_132 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U1 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 
+ TSMC_261 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 TSMC_243 
+ TSMC_244 TSMC_245 TSMC_36 TSMC_68 TSMC_100 TSMC_132 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D2 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 TSMC_283 TSMC_284 
+ TSMC_285 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 
+ TSMC_268 TSMC_269 TSMC_37 TSMC_69 TSMC_101 TSMC_133 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U2 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 TSMC_291 TSMC_292 
+ TSMC_293 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 TSMC_275 
+ TSMC_276 TSMC_277 TSMC_37 TSMC_69 TSMC_101 TSMC_133 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D3 TSMC_310 TSMC_311 TSMC_312 TSMC_313 TSMC_314 TSMC_315 TSMC_316 
+ TSMC_317 TSMC_294 TSMC_295 TSMC_296 TSMC_297 TSMC_298 TSMC_299 
+ TSMC_300 TSMC_301 TSMC_38 TSMC_70 TSMC_102 TSMC_134 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U3 TSMC_318 TSMC_319 TSMC_320 TSMC_321 TSMC_322 TSMC_323 TSMC_324 
+ TSMC_325 TSMC_302 TSMC_303 TSMC_304 TSMC_305 TSMC_306 TSMC_307 
+ TSMC_308 TSMC_309 TSMC_38 TSMC_70 TSMC_102 TSMC_134 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D4 TSMC_342 TSMC_343 TSMC_344 TSMC_345 TSMC_346 TSMC_347 TSMC_348 
+ TSMC_349 TSMC_326 TSMC_327 TSMC_328 TSMC_329 TSMC_330 TSMC_331 
+ TSMC_332 TSMC_333 TSMC_39 TSMC_71 TSMC_103 TSMC_135 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U4 TSMC_350 TSMC_351 TSMC_352 TSMC_353 TSMC_354 TSMC_355 TSMC_356 
+ TSMC_357 TSMC_334 TSMC_335 TSMC_336 TSMC_337 TSMC_338 TSMC_339 
+ TSMC_340 TSMC_341 TSMC_39 TSMC_71 TSMC_103 TSMC_135 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D5 TSMC_374 TSMC_375 TSMC_376 TSMC_377 TSMC_378 TSMC_379 TSMC_380 
+ TSMC_381 TSMC_358 TSMC_359 TSMC_360 TSMC_361 TSMC_362 TSMC_363 
+ TSMC_364 TSMC_365 TSMC_40 TSMC_72 TSMC_104 TSMC_136 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U5 TSMC_382 TSMC_383 TSMC_384 TSMC_385 TSMC_386 TSMC_387 TSMC_388 
+ TSMC_389 TSMC_366 TSMC_367 TSMC_368 TSMC_369 TSMC_370 TSMC_371 
+ TSMC_372 TSMC_373 TSMC_40 TSMC_72 TSMC_104 TSMC_136 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D6 TSMC_406 TSMC_407 TSMC_408 TSMC_409 TSMC_410 TSMC_411 TSMC_412 
+ TSMC_413 TSMC_390 TSMC_391 TSMC_392 TSMC_393 TSMC_394 TSMC_395 
+ TSMC_396 TSMC_397 TSMC_41 TSMC_73 TSMC_105 TSMC_137 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U6 TSMC_414 TSMC_415 TSMC_416 TSMC_417 TSMC_418 TSMC_419 TSMC_420 
+ TSMC_421 TSMC_398 TSMC_399 TSMC_400 TSMC_401 TSMC_402 TSMC_403 
+ TSMC_404 TSMC_405 TSMC_41 TSMC_73 TSMC_105 TSMC_137 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D7 TSMC_438 TSMC_439 TSMC_440 TSMC_441 TSMC_442 TSMC_443 TSMC_444 
+ TSMC_445 TSMC_422 TSMC_423 TSMC_424 TSMC_425 TSMC_426 TSMC_427 
+ TSMC_428 TSMC_429 TSMC_42 TSMC_74 TSMC_106 TSMC_138 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U7 TSMC_446 TSMC_447 TSMC_448 TSMC_449 TSMC_450 TSMC_451 TSMC_452 
+ TSMC_453 TSMC_430 TSMC_431 TSMC_432 TSMC_433 TSMC_434 TSMC_435 
+ TSMC_436 TSMC_437 TSMC_42 TSMC_74 TSMC_106 TSMC_138 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D8 TSMC_470 TSMC_471 TSMC_472 TSMC_473 TSMC_474 TSMC_475 TSMC_476 
+ TSMC_477 TSMC_454 TSMC_455 TSMC_456 TSMC_457 TSMC_458 TSMC_459 
+ TSMC_460 TSMC_461 TSMC_43 TSMC_75 TSMC_107 TSMC_139 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U8 TSMC_478 TSMC_479 TSMC_480 TSMC_481 TSMC_482 TSMC_483 TSMC_484 
+ TSMC_485 TSMC_462 TSMC_463 TSMC_464 TSMC_465 TSMC_466 TSMC_467 
+ TSMC_468 TSMC_469 TSMC_43 TSMC_75 TSMC_107 TSMC_139 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D9 TSMC_502 TSMC_503 TSMC_504 TSMC_505 TSMC_506 TSMC_507 TSMC_508 
+ TSMC_509 TSMC_486 TSMC_487 TSMC_488 TSMC_489 TSMC_490 TSMC_491 
+ TSMC_492 TSMC_493 TSMC_44 TSMC_76 TSMC_108 TSMC_140 VDDAI VDDI VSSI TSMC_1248 
+ TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 TSMC_1293 
+ TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 TSMC_1325 
+ TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 TSMC_1357 
+ TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 TSMC_1401 
+ TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 TSMC_1420 
+ TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 TSMC_1464 
+ TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 TSMC_1483 
+ TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U9 TSMC_510 TSMC_511 TSMC_512 TSMC_513 TSMC_514 TSMC_515 TSMC_516 
+ TSMC_517 TSMC_494 TSMC_495 TSMC_496 TSMC_497 TSMC_498 TSMC_499 
+ TSMC_500 TSMC_501 TSMC_44 TSMC_76 TSMC_108 TSMC_140 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 TSMC_1552 
+ TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 TSMC_1615 
+ TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 TSMC_1678 
+ TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 TSMC_1741 
+ TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D10 TSMC_534 TSMC_535 TSMC_536 TSMC_537 TSMC_538 TSMC_539 
+ TSMC_540 TSMC_541 TSMC_518 TSMC_519 TSMC_520 TSMC_521 TSMC_522 
+ TSMC_523 TSMC_524 TSMC_525 TSMC_45 TSMC_77 TSMC_109 TSMC_141 VDDAI VDDI VSSI 
+ TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U10 TSMC_542 TSMC_543 TSMC_544 TSMC_545 TSMC_546 TSMC_547 
+ TSMC_548 TSMC_549 TSMC_526 TSMC_527 TSMC_528 TSMC_529 TSMC_530 
+ TSMC_531 TSMC_532 TSMC_533 TSMC_45 TSMC_77 TSMC_109 TSMC_141 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 
+ TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 
+ TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 
+ TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 
+ TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 
+ TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 
+ TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 
+ TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 
+ TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 
+ TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D11 TSMC_566 TSMC_567 TSMC_568 TSMC_569 TSMC_570 TSMC_571 
+ TSMC_572 TSMC_573 TSMC_550 TSMC_551 TSMC_552 TSMC_553 TSMC_554 
+ TSMC_555 TSMC_556 TSMC_557 TSMC_46 TSMC_78 TSMC_110 TSMC_142 VDDAI VDDI VSSI 
+ TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 
+ TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 
+ TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 
+ TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 
+ TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U11 TSMC_574 TSMC_575 TSMC_576 TSMC_577 TSMC_578 TSMC_579 
+ TSMC_580 TSMC_581 TSMC_558 TSMC_559 TSMC_560 TSMC_561 TSMC_562 
+ TSMC_563 TSMC_564 TSMC_565 TSMC_46 TSMC_78 TSMC_110 TSMC_142 VDDAI VDDI VSSI 
+ TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 
+ TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 
+ TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 
+ TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 
+ TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 
+ TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 
+ TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 
+ TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 
+ TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 
+ TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 
+ TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D12 TSMC_598 TSMC_599 TSMC_600 TSMC_601 TSMC_602 TSMC_603 
+ TSMC_604 TSMC_605 TSMC_582 TSMC_583 TSMC_584 TSMC_585 TSMC_586 
+ TSMC_587 TSMC_588 TSMC_589 TSMC_47 TSMC_79 TSMC_111 TSMC_143 VDDAI VDDI 
+ VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 TSMC_1254 
+ TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 TSMC_1260 
+ TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 TSMC_1267 
+ TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 TSMC_1273 
+ TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 TSMC_1279 TSMC_1280 
+ TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 TSMC_1286 
+ TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 TSMC_1292 
+ TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 TSMC_1299 
+ TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 TSMC_1305 
+ TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 TSMC_1311 TSMC_1312 
+ TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 TSMC_1318 
+ TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 TSMC_1324 
+ TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 TSMC_1331 
+ TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 TSMC_1337 
+ TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 TSMC_1344 
+ TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 TSMC_1350 
+ TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 TSMC_1356 
+ TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 TSMC_1363 
+ TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 TSMC_1369 
+ TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 TSMC_1375 
+ TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 TSMC_1381 TSMC_1382 
+ TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 TSMC_1388 
+ TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 TSMC_1394 
+ TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 TSMC_1400 
+ TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 TSMC_1407 
+ TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 TSMC_1413 
+ TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 TSMC_1419 
+ TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 TSMC_1426 
+ TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 TSMC_1432 
+ TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 TSMC_1438 
+ TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 TSMC_1444 TSMC_1445 
+ TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 TSMC_1451 
+ TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 TSMC_1457 
+ TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 TSMC_1463 
+ TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 TSMC_1470 
+ TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 TSMC_1476 
+ TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 TSMC_1482 
+ TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 TSMC_1489 
+ TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 TSMC_1495 
+ TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 TSMC_1501 
+ TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U12 TSMC_606 TSMC_607 TSMC_608 TSMC_609 TSMC_610 TSMC_611 
+ TSMC_612 TSMC_613 TSMC_590 TSMC_591 TSMC_592 TSMC_593 TSMC_594 
+ TSMC_595 TSMC_596 TSMC_597 TSMC_47 TSMC_79 TSMC_111 TSMC_143 VDDAI VDDI 
+ VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 TSMC_1513 TSMC_1514 
+ TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 TSMC_1520 
+ TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 TSMC_1526 
+ TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 TSMC_1532 TSMC_1533 
+ TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 TSMC_1539 
+ TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 TSMC_1545 
+ TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 TSMC_1551 
+ TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 TSMC_1558 
+ TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 TSMC_1564 
+ TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 TSMC_1570 
+ TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 TSMC_1576 TSMC_1577 
+ TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 TSMC_1583 
+ TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 TSMC_1589 
+ TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 TSMC_1595 TSMC_1596 
+ TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 TSMC_1602 
+ TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 TSMC_1608 
+ TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 TSMC_1614 
+ TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 TSMC_1621 
+ TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 TSMC_1627 
+ TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 TSMC_1633 
+ TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 TSMC_1639 TSMC_1640 
+ TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 TSMC_1646 
+ TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 TSMC_1652 
+ TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 TSMC_1658 TSMC_1659 
+ TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 TSMC_1665 
+ TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 TSMC_1671 
+ TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 TSMC_1677 
+ TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 TSMC_1684 
+ TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 TSMC_1690 
+ TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 TSMC_1696 
+ TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 TSMC_1702 TSMC_1703 
+ TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 TSMC_1709 
+ TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 TSMC_1715 
+ TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 TSMC_1721 TSMC_1722 
+ TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 TSMC_1728 
+ TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 TSMC_1734 
+ TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 TSMC_1740 
+ TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 TSMC_1747 
+ TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 TSMC_1753 
+ TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 TSMC_1759 
+ TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D13 TSMC_630 TSMC_631 TSMC_632 TSMC_633 TSMC_634 TSMC_635 
+ TSMC_636 TSMC_637 TSMC_614 TSMC_615 TSMC_616 TSMC_617 TSMC_618 
+ TSMC_619 TSMC_620 TSMC_621 TSMC_48 TSMC_80 TSMC_112 TSMC_144 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U13 TSMC_638 TSMC_639 TSMC_640 TSMC_641 TSMC_642 TSMC_643 
+ TSMC_644 TSMC_645 TSMC_622 TSMC_623 TSMC_624 TSMC_625 TSMC_626 
+ TSMC_627 TSMC_628 TSMC_629 TSMC_48 TSMC_80 TSMC_112 TSMC_144 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D14 TSMC_662 TSMC_663 TSMC_664 TSMC_665 TSMC_666 TSMC_667 
+ TSMC_668 TSMC_669 TSMC_646 TSMC_647 TSMC_648 TSMC_649 TSMC_650 
+ TSMC_651 TSMC_652 TSMC_653 TSMC_49 TSMC_81 TSMC_113 TSMC_145 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U14 TSMC_670 TSMC_671 TSMC_672 TSMC_673 TSMC_674 TSMC_675 
+ TSMC_676 TSMC_677 TSMC_654 TSMC_655 TSMC_656 TSMC_657 TSMC_658 
+ TSMC_659 TSMC_660 TSMC_661 TSMC_49 TSMC_81 TSMC_113 TSMC_145 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D15 TSMC_694 TSMC_695 TSMC_696 TSMC_697 TSMC_698 TSMC_699 
+ TSMC_700 TSMC_701 TSMC_678 TSMC_679 TSMC_680 TSMC_681 TSMC_682 
+ TSMC_683 TSMC_684 TSMC_685 TSMC_50 TSMC_82 TSMC_114 TSMC_146 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U15 TSMC_702 TSMC_703 TSMC_704 TSMC_705 TSMC_706 TSMC_707 
+ TSMC_708 TSMC_709 TSMC_686 TSMC_687 TSMC_688 TSMC_689 TSMC_690 
+ TSMC_691 TSMC_692 TSMC_693 TSMC_50 TSMC_82 TSMC_114 TSMC_146 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D16 TSMC_726 TSMC_727 TSMC_728 TSMC_729 TSMC_730 TSMC_731 
+ TSMC_732 TSMC_733 TSMC_710 TSMC_711 TSMC_712 TSMC_713 TSMC_714 
+ TSMC_715 TSMC_716 TSMC_717 TSMC_51 TSMC_83 TSMC_115 TSMC_147 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U16 TSMC_734 TSMC_735 TSMC_736 TSMC_737 TSMC_738 TSMC_739 
+ TSMC_740 TSMC_741 TSMC_718 TSMC_719 TSMC_720 TSMC_721 TSMC_722 
+ TSMC_723 TSMC_724 TSMC_725 TSMC_51 TSMC_83 TSMC_115 TSMC_147 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D17 TSMC_758 TSMC_759 TSMC_760 TSMC_761 TSMC_762 TSMC_763 
+ TSMC_764 TSMC_765 TSMC_742 TSMC_743 TSMC_744 TSMC_745 TSMC_746 
+ TSMC_747 TSMC_748 TSMC_749 TSMC_52 TSMC_84 TSMC_116 TSMC_148 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U17 TSMC_766 TSMC_767 TSMC_768 TSMC_769 TSMC_770 TSMC_771 
+ TSMC_772 TSMC_773 TSMC_750 TSMC_751 TSMC_752 TSMC_753 TSMC_754 
+ TSMC_755 TSMC_756 TSMC_757 TSMC_52 TSMC_84 TSMC_116 TSMC_148 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D18 TSMC_790 TSMC_791 TSMC_792 TSMC_793 TSMC_794 TSMC_795 
+ TSMC_796 TSMC_797 TSMC_774 TSMC_775 TSMC_776 TSMC_777 TSMC_778 
+ TSMC_779 TSMC_780 TSMC_781 TSMC_53 TSMC_85 TSMC_117 TSMC_149 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U18 TSMC_798 TSMC_799 TSMC_800 TSMC_801 TSMC_802 TSMC_803 
+ TSMC_804 TSMC_805 TSMC_782 TSMC_783 TSMC_784 TSMC_785 TSMC_786 
+ TSMC_787 TSMC_788 TSMC_789 TSMC_53 TSMC_85 TSMC_117 TSMC_149 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D19 TSMC_822 TSMC_823 TSMC_824 TSMC_825 TSMC_826 TSMC_827 
+ TSMC_828 TSMC_829 TSMC_806 TSMC_807 TSMC_808 TSMC_809 TSMC_810 
+ TSMC_811 TSMC_812 TSMC_813 TSMC_54 TSMC_86 TSMC_118 TSMC_150 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U19 TSMC_830 TSMC_831 TSMC_832 TSMC_833 TSMC_834 TSMC_835 
+ TSMC_836 TSMC_837 TSMC_814 TSMC_815 TSMC_816 TSMC_817 TSMC_818 
+ TSMC_819 TSMC_820 TSMC_821 TSMC_54 TSMC_86 TSMC_118 TSMC_150 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D20 TSMC_854 TSMC_855 TSMC_856 TSMC_857 TSMC_858 TSMC_859 
+ TSMC_860 TSMC_861 TSMC_838 TSMC_839 TSMC_840 TSMC_841 TSMC_842 
+ TSMC_843 TSMC_844 TSMC_845 TSMC_55 TSMC_87 TSMC_119 TSMC_151 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U20 TSMC_862 TSMC_863 TSMC_864 TSMC_865 TSMC_866 TSMC_867 
+ TSMC_868 TSMC_869 TSMC_846 TSMC_847 TSMC_848 TSMC_849 TSMC_850 
+ TSMC_851 TSMC_852 TSMC_853 TSMC_55 TSMC_87 TSMC_119 TSMC_151 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D21 TSMC_886 TSMC_887 TSMC_888 TSMC_889 TSMC_890 TSMC_891 
+ TSMC_892 TSMC_893 TSMC_870 TSMC_871 TSMC_872 TSMC_873 TSMC_874 
+ TSMC_875 TSMC_876 TSMC_877 TSMC_56 TSMC_88 TSMC_120 TSMC_152 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U21 TSMC_894 TSMC_895 TSMC_896 TSMC_897 TSMC_898 TSMC_899 
+ TSMC_900 TSMC_901 TSMC_878 TSMC_879 TSMC_880 TSMC_881 TSMC_882 
+ TSMC_883 TSMC_884 TSMC_885 TSMC_56 TSMC_88 TSMC_120 TSMC_152 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D22 TSMC_918 TSMC_919 TSMC_920 TSMC_921 TSMC_922 TSMC_923 
+ TSMC_924 TSMC_925 TSMC_902 TSMC_903 TSMC_904 TSMC_905 TSMC_906 
+ TSMC_907 TSMC_908 TSMC_909 TSMC_57 TSMC_89 TSMC_121 TSMC_153 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U22 TSMC_926 TSMC_927 TSMC_928 TSMC_929 TSMC_930 TSMC_931 
+ TSMC_932 TSMC_933 TSMC_910 TSMC_911 TSMC_912 TSMC_913 TSMC_914 
+ TSMC_915 TSMC_916 TSMC_917 TSMC_57 TSMC_89 TSMC_121 TSMC_153 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D23 TSMC_950 TSMC_951 TSMC_952 TSMC_953 TSMC_954 TSMC_955 
+ TSMC_956 TSMC_957 TSMC_934 TSMC_935 TSMC_936 TSMC_937 TSMC_938 
+ TSMC_939 TSMC_940 TSMC_941 TSMC_58 TSMC_90 TSMC_122 TSMC_154 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U23 TSMC_958 TSMC_959 TSMC_960 TSMC_961 TSMC_962 TSMC_963 
+ TSMC_964 TSMC_965 TSMC_942 TSMC_943 TSMC_944 TSMC_945 TSMC_946 
+ TSMC_947 TSMC_948 TSMC_949 TSMC_58 TSMC_90 TSMC_122 TSMC_154 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D24 TSMC_982 TSMC_983 TSMC_984 TSMC_985 TSMC_986 TSMC_987 
+ TSMC_988 TSMC_989 TSMC_966 TSMC_967 TSMC_968 TSMC_969 TSMC_970 
+ TSMC_971 TSMC_972 TSMC_973 TSMC_59 TSMC_91 TSMC_123 TSMC_155 VDDAI 
+ VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U24 TSMC_990 TSMC_991 TSMC_992 TSMC_993 TSMC_994 TSMC_995 
+ TSMC_996 TSMC_997 TSMC_974 TSMC_975 TSMC_976 TSMC_977 TSMC_978 
+ TSMC_979 TSMC_980 TSMC_981 TSMC_59 TSMC_91 TSMC_123 TSMC_155 VDDAI 
+ VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 TSMC_1519 
+ TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 TSMC_1525 
+ TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 TSMC_1531 
+ TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 TSMC_1538 
+ TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 TSMC_1544 
+ TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 TSMC_1550 
+ TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 TSMC_1557 
+ TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 TSMC_1563 
+ TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 TSMC_1569 
+ TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 TSMC_1582 
+ TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 TSMC_1588 
+ TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 TSMC_1594 
+ TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 TSMC_1601 
+ TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 TSMC_1607 
+ TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 TSMC_1613 
+ TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 TSMC_1620 
+ TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 TSMC_1626 
+ TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 TSMC_1632 
+ TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 TSMC_1645 
+ TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 TSMC_1651 
+ TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 TSMC_1657 
+ TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 TSMC_1664 
+ TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 TSMC_1670 
+ TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 TSMC_1676 
+ TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 TSMC_1683 
+ TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 TSMC_1689 
+ TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 TSMC_1695 
+ TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 TSMC_1708 
+ TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 TSMC_1714 
+ TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 TSMC_1720 
+ TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 TSMC_1727 
+ TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 TSMC_1733 
+ TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 TSMC_1739 
+ TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 TSMC_1746 
+ TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 TSMC_1752 
+ TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 TSMC_1758 
+ TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D25 TSMC_1014 TSMC_1015 TSMC_1016 TSMC_1017 TSMC_1018 TSMC_1019 
+ TSMC_1020 TSMC_1021 TSMC_998 TSMC_999 TSMC_1000 TSMC_1001 TSMC_1002 
+ TSMC_1003 TSMC_1004 TSMC_1005 TSMC_60 TSMC_92 TSMC_124 TSMC_156 
+ VDDAI VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 TSMC_1253 
+ TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 TSMC_1259 
+ TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 TSMC_1266 
+ TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 TSMC_1272 
+ TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 TSMC_1278 
+ TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 TSMC_1285 
+ TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 TSMC_1291 
+ TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 TSMC_1298 
+ TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 TSMC_1304 
+ TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 TSMC_1317 
+ TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 TSMC_1323 
+ TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 TSMC_1330 
+ TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 TSMC_1336 
+ TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 TSMC_1343 
+ TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 TSMC_1349 
+ TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 TSMC_1355 
+ TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 TSMC_1362 
+ TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 TSMC_1368 
+ TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 TSMC_1374 
+ TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 TSMC_1387 
+ TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 TSMC_1393 
+ TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 TSMC_1399 
+ TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 TSMC_1406 
+ TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 TSMC_1412 
+ TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 TSMC_1418 
+ TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 TSMC_1425 
+ TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 TSMC_1431 
+ TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 TSMC_1437 
+ TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 TSMC_1450 
+ TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 TSMC_1456 
+ TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 TSMC_1462 
+ TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 TSMC_1469 
+ TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 TSMC_1475 
+ TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 TSMC_1481 
+ TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 TSMC_1488 
+ TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 TSMC_1494 
+ TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 TSMC_1500 
+ TSMC_1501 TSMC_1502 TSMC_1503 S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U25 TSMC_1022 TSMC_1023 TSMC_1024 TSMC_1025 TSMC_1026 TSMC_1027 
+ TSMC_1028 TSMC_1029 TSMC_1006 TSMC_1007 TSMC_1008 TSMC_1009 
+ TSMC_1010 TSMC_1011 TSMC_1012 TSMC_1013 TSMC_60 TSMC_92 TSMC_124 
+ TSMC_156 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D26 TSMC_1046 TSMC_1047 TSMC_1048 TSMC_1049 TSMC_1050 TSMC_1051 
+ TSMC_1052 TSMC_1053 TSMC_1030 TSMC_1031 TSMC_1032 TSMC_1033 
+ TSMC_1034 TSMC_1035 TSMC_1036 TSMC_1037 TSMC_61 TSMC_93 TSMC_125 
+ TSMC_157 VDDAI VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 
+ TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 
+ TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 
+ TSMC_1272 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 
+ TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 
+ TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 
+ TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 
+ TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 
+ TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 
+ TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 
+ TSMC_1336 TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 
+ TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 
+ TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 
+ TSMC_1368 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 
+ TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 
+ TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 
+ TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 
+ TSMC_1412 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 
+ TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 
+ TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 
+ TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 
+ TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 
+ TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 
+ TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 
+ TSMC_1488 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 
+ TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U26 TSMC_1054 TSMC_1055 TSMC_1056 TSMC_1057 TSMC_1058 TSMC_1059 
+ TSMC_1060 TSMC_1061 TSMC_1038 TSMC_1039 TSMC_1040 TSMC_1041 
+ TSMC_1042 TSMC_1043 TSMC_1044 TSMC_1045 TSMC_61 TSMC_93 TSMC_125 
+ TSMC_157 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D27 TSMC_1078 TSMC_1079 TSMC_1080 TSMC_1081 TSMC_1082 TSMC_1083 
+ TSMC_1084 TSMC_1085 TSMC_1062 TSMC_1063 TSMC_1064 TSMC_1065 
+ TSMC_1066 TSMC_1067 TSMC_1068 TSMC_1069 TSMC_62 TSMC_94 TSMC_126 
+ TSMC_158 VDDAI VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 
+ TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 
+ TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 
+ TSMC_1272 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 
+ TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 
+ TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 
+ TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 
+ TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 
+ TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 
+ TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 
+ TSMC_1336 TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 
+ TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 
+ TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 
+ TSMC_1368 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 
+ TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 
+ TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 
+ TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 
+ TSMC_1412 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 
+ TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 
+ TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 
+ TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 
+ TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 
+ TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 
+ TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 
+ TSMC_1488 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 
+ TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U27 TSMC_1086 TSMC_1087 TSMC_1088 TSMC_1089 TSMC_1090 TSMC_1091 
+ TSMC_1092 TSMC_1093 TSMC_1070 TSMC_1071 TSMC_1072 TSMC_1073 
+ TSMC_1074 TSMC_1075 TSMC_1076 TSMC_1077 TSMC_62 TSMC_94 TSMC_126 
+ TSMC_158 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D28 TSMC_1110 TSMC_1111 TSMC_1112 TSMC_1113 TSMC_1114 TSMC_1115 
+ TSMC_1116 TSMC_1117 TSMC_1094 TSMC_1095 TSMC_1096 TSMC_1097 
+ TSMC_1098 TSMC_1099 TSMC_1100 TSMC_1101 TSMC_63 TSMC_95 TSMC_127 
+ TSMC_159 VDDAI VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 
+ TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 
+ TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 
+ TSMC_1272 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 
+ TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 
+ TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 
+ TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 
+ TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 
+ TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 
+ TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 
+ TSMC_1336 TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 
+ TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 
+ TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 
+ TSMC_1368 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 
+ TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 
+ TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 
+ TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 
+ TSMC_1412 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 
+ TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 
+ TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 
+ TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 
+ TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 
+ TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 
+ TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 
+ TSMC_1488 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 
+ TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U28 TSMC_1118 TSMC_1119 TSMC_1120 TSMC_1121 TSMC_1122 TSMC_1123 
+ TSMC_1124 TSMC_1125 TSMC_1102 TSMC_1103 TSMC_1104 TSMC_1105 
+ TSMC_1106 TSMC_1107 TSMC_1108 TSMC_1109 TSMC_63 TSMC_95 TSMC_127 
+ TSMC_159 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D29 TSMC_1142 TSMC_1143 TSMC_1144 TSMC_1145 TSMC_1146 TSMC_1147 
+ TSMC_1148 TSMC_1149 TSMC_1126 TSMC_1127 TSMC_1128 TSMC_1129 
+ TSMC_1130 TSMC_1131 TSMC_1132 TSMC_1133 TSMC_64 TSMC_96 TSMC_128 
+ TSMC_160 VDDAI VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 
+ TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 
+ TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 
+ TSMC_1272 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 
+ TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 
+ TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 
+ TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 
+ TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 
+ TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 
+ TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 
+ TSMC_1336 TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 
+ TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 
+ TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 
+ TSMC_1368 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 
+ TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 
+ TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 
+ TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 
+ TSMC_1412 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 
+ TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 
+ TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 
+ TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 
+ TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 
+ TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 
+ TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 
+ TSMC_1488 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 
+ TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U29 TSMC_1150 TSMC_1151 TSMC_1152 TSMC_1153 TSMC_1154 TSMC_1155 
+ TSMC_1156 TSMC_1157 TSMC_1134 TSMC_1135 TSMC_1136 TSMC_1137 
+ TSMC_1138 TSMC_1139 TSMC_1140 TSMC_1141 TSMC_64 TSMC_96 TSMC_128 
+ TSMC_160 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D30 TSMC_1174 TSMC_1175 TSMC_1176 TSMC_1177 TSMC_1178 TSMC_1179 
+ TSMC_1180 TSMC_1181 TSMC_1158 TSMC_1159 TSMC_1160 TSMC_1161 
+ TSMC_1162 TSMC_1163 TSMC_1164 TSMC_1165 TSMC_65 TSMC_97 TSMC_129 
+ TSMC_161 VDDAI VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 
+ TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 
+ TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 
+ TSMC_1272 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 
+ TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 
+ TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 
+ TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 
+ TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 
+ TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 
+ TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 
+ TSMC_1336 TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 
+ TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 
+ TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 
+ TSMC_1368 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 
+ TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 
+ TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 
+ TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 
+ TSMC_1412 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 
+ TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 
+ TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 
+ TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 
+ TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 
+ TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 
+ TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 
+ TSMC_1488 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 
+ TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U30 TSMC_1182 TSMC_1183 TSMC_1184 TSMC_1185 TSMC_1186 TSMC_1187 
+ TSMC_1188 TSMC_1189 TSMC_1166 TSMC_1167 TSMC_1168 TSMC_1169 
+ TSMC_1170 TSMC_1171 TSMC_1172 TSMC_1173 TSMC_65 TSMC_97 TSMC_129 
+ TSMC_161 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_D31 TSMC_1206 TSMC_1207 TSMC_1208 TSMC_1209 TSMC_1210 TSMC_1211 
+ TSMC_1212 TSMC_1213 TSMC_1190 TSMC_1191 TSMC_1192 TSMC_1193 
+ TSMC_1194 TSMC_1195 TSMC_1196 TSMC_1197 TSMC_66 TSMC_98 TSMC_130 
+ TSMC_162 VDDAI VDDI VSSI TSMC_1248 TSMC_1249 TSMC_1250 TSMC_1251 TSMC_1252 
+ TSMC_1253 TSMC_1254 TSMC_1255 TSMC_1256 TSMC_1257 TSMC_1258 
+ TSMC_1259 TSMC_1260 TSMC_1261 TSMC_1262 TSMC_1263 TSMC_1264 TSMC_1265 
+ TSMC_1266 TSMC_1267 TSMC_1268 TSMC_1269 TSMC_1270 TSMC_1271 
+ TSMC_1272 TSMC_1273 TSMC_1274 TSMC_1275 TSMC_1276 TSMC_1277 
+ TSMC_1278 TSMC_1279 TSMC_1280 TSMC_1281 TSMC_1282 TSMC_1283 TSMC_1284 
+ TSMC_1285 TSMC_1286 TSMC_1287 TSMC_1288 TSMC_1289 TSMC_1290 
+ TSMC_1291 TSMC_1292 TSMC_1293 TSMC_1294 TSMC_1295 TSMC_1296 TSMC_1297 
+ TSMC_1298 TSMC_1299 TSMC_1300 TSMC_1301 TSMC_1302 TSMC_1303 
+ TSMC_1304 TSMC_1305 TSMC_1306 TSMC_1307 TSMC_1308 TSMC_1309 TSMC_1310 
+ TSMC_1311 TSMC_1312 TSMC_1313 TSMC_1314 TSMC_1315 TSMC_1316 
+ TSMC_1317 TSMC_1318 TSMC_1319 TSMC_1320 TSMC_1321 TSMC_1322 
+ TSMC_1323 TSMC_1324 TSMC_1325 TSMC_1326 TSMC_1327 TSMC_1328 TSMC_1329 
+ TSMC_1330 TSMC_1331 TSMC_1332 TSMC_1333 TSMC_1334 TSMC_1335 
+ TSMC_1336 TSMC_1337 TSMC_1338 TSMC_1339 TSMC_1340 TSMC_1341 TSMC_1342 
+ TSMC_1343 TSMC_1344 TSMC_1345 TSMC_1346 TSMC_1347 TSMC_1348 
+ TSMC_1349 TSMC_1350 TSMC_1351 TSMC_1352 TSMC_1353 TSMC_1354 
+ TSMC_1355 TSMC_1356 TSMC_1357 TSMC_1358 TSMC_1359 TSMC_1360 TSMC_1361 
+ TSMC_1362 TSMC_1363 TSMC_1364 TSMC_1365 TSMC_1366 TSMC_1367 
+ TSMC_1368 TSMC_1369 TSMC_1370 TSMC_1371 TSMC_1372 TSMC_1373 
+ TSMC_1374 TSMC_1375 TSMC_1376 TSMC_1377 TSMC_1378 TSMC_1379 TSMC_1380 
+ TSMC_1381 TSMC_1382 TSMC_1383 TSMC_1384 TSMC_1385 TSMC_1386 
+ TSMC_1387 TSMC_1388 TSMC_1389 TSMC_1390 TSMC_1391 TSMC_1392 
+ TSMC_1393 TSMC_1394 TSMC_1395 TSMC_1396 TSMC_1397 TSMC_1398 
+ TSMC_1399 TSMC_1400 TSMC_1401 TSMC_1402 TSMC_1403 TSMC_1404 TSMC_1405 
+ TSMC_1406 TSMC_1407 TSMC_1408 TSMC_1409 TSMC_1410 TSMC_1411 
+ TSMC_1412 TSMC_1413 TSMC_1414 TSMC_1415 TSMC_1416 TSMC_1417 
+ TSMC_1418 TSMC_1419 TSMC_1420 TSMC_1421 TSMC_1422 TSMC_1423 TSMC_1424 
+ TSMC_1425 TSMC_1426 TSMC_1427 TSMC_1428 TSMC_1429 TSMC_1430 
+ TSMC_1431 TSMC_1432 TSMC_1433 TSMC_1434 TSMC_1435 TSMC_1436 
+ TSMC_1437 TSMC_1438 TSMC_1439 TSMC_1440 TSMC_1441 TSMC_1442 TSMC_1443 
+ TSMC_1444 TSMC_1445 TSMC_1446 TSMC_1447 TSMC_1448 TSMC_1449 
+ TSMC_1450 TSMC_1451 TSMC_1452 TSMC_1453 TSMC_1454 TSMC_1455 
+ TSMC_1456 TSMC_1457 TSMC_1458 TSMC_1459 TSMC_1460 TSMC_1461 
+ TSMC_1462 TSMC_1463 TSMC_1464 TSMC_1465 TSMC_1466 TSMC_1467 TSMC_1468 
+ TSMC_1469 TSMC_1470 TSMC_1471 TSMC_1472 TSMC_1473 TSMC_1474 
+ TSMC_1475 TSMC_1476 TSMC_1477 TSMC_1478 TSMC_1479 TSMC_1480 
+ TSMC_1481 TSMC_1482 TSMC_1483 TSMC_1484 TSMC_1485 TSMC_1486 TSMC_1487 
+ TSMC_1488 TSMC_1489 TSMC_1490 TSMC_1491 TSMC_1492 TSMC_1493 
+ TSMC_1494 TSMC_1495 TSMC_1496 TSMC_1497 TSMC_1498 TSMC_1499 
+ TSMC_1500 TSMC_1501 TSMC_1502 TSMC_1503 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
XMCB_U31 TSMC_1214 TSMC_1215 TSMC_1216 TSMC_1217 TSMC_1218 TSMC_1219 
+ TSMC_1220 TSMC_1221 TSMC_1198 TSMC_1199 TSMC_1200 TSMC_1201 
+ TSMC_1202 TSMC_1203 TSMC_1204 TSMC_1205 TSMC_66 TSMC_98 TSMC_130 
+ TSMC_162 VDDAI VDDI VSSI TSMC_1508 TSMC_1509 TSMC_1510 TSMC_1511 TSMC_1512 
+ TSMC_1513 TSMC_1514 TSMC_1515 TSMC_1516 TSMC_1517 TSMC_1518 
+ TSMC_1519 TSMC_1520 TSMC_1521 TSMC_1522 TSMC_1523 TSMC_1524 
+ TSMC_1525 TSMC_1526 TSMC_1527 TSMC_1528 TSMC_1529 TSMC_1530 
+ TSMC_1531 TSMC_1532 TSMC_1533 TSMC_1534 TSMC_1535 TSMC_1536 TSMC_1537 
+ TSMC_1538 TSMC_1539 TSMC_1540 TSMC_1541 TSMC_1542 TSMC_1543 
+ TSMC_1544 TSMC_1545 TSMC_1546 TSMC_1547 TSMC_1548 TSMC_1549 
+ TSMC_1550 TSMC_1551 TSMC_1552 TSMC_1553 TSMC_1554 TSMC_1555 TSMC_1556 
+ TSMC_1557 TSMC_1558 TSMC_1559 TSMC_1560 TSMC_1561 TSMC_1562 
+ TSMC_1563 TSMC_1564 TSMC_1565 TSMC_1566 TSMC_1567 TSMC_1568 
+ TSMC_1569 TSMC_1570 TSMC_1571 TSMC_1572 TSMC_1573 TSMC_1574 TSMC_1575 
+ TSMC_1576 TSMC_1577 TSMC_1578 TSMC_1579 TSMC_1580 TSMC_1581 
+ TSMC_1582 TSMC_1583 TSMC_1584 TSMC_1585 TSMC_1586 TSMC_1587 
+ TSMC_1588 TSMC_1589 TSMC_1590 TSMC_1591 TSMC_1592 TSMC_1593 
+ TSMC_1594 TSMC_1595 TSMC_1596 TSMC_1597 TSMC_1598 TSMC_1599 TSMC_1600 
+ TSMC_1601 TSMC_1602 TSMC_1603 TSMC_1604 TSMC_1605 TSMC_1606 
+ TSMC_1607 TSMC_1608 TSMC_1609 TSMC_1610 TSMC_1611 TSMC_1612 
+ TSMC_1613 TSMC_1614 TSMC_1615 TSMC_1616 TSMC_1617 TSMC_1618 TSMC_1619 
+ TSMC_1620 TSMC_1621 TSMC_1622 TSMC_1623 TSMC_1624 TSMC_1625 
+ TSMC_1626 TSMC_1627 TSMC_1628 TSMC_1629 TSMC_1630 TSMC_1631 
+ TSMC_1632 TSMC_1633 TSMC_1634 TSMC_1635 TSMC_1636 TSMC_1637 TSMC_1638 
+ TSMC_1639 TSMC_1640 TSMC_1641 TSMC_1642 TSMC_1643 TSMC_1644 
+ TSMC_1645 TSMC_1646 TSMC_1647 TSMC_1648 TSMC_1649 TSMC_1650 
+ TSMC_1651 TSMC_1652 TSMC_1653 TSMC_1654 TSMC_1655 TSMC_1656 
+ TSMC_1657 TSMC_1658 TSMC_1659 TSMC_1660 TSMC_1661 TSMC_1662 TSMC_1663 
+ TSMC_1664 TSMC_1665 TSMC_1666 TSMC_1667 TSMC_1668 TSMC_1669 
+ TSMC_1670 TSMC_1671 TSMC_1672 TSMC_1673 TSMC_1674 TSMC_1675 
+ TSMC_1676 TSMC_1677 TSMC_1678 TSMC_1679 TSMC_1680 TSMC_1681 TSMC_1682 
+ TSMC_1683 TSMC_1684 TSMC_1685 TSMC_1686 TSMC_1687 TSMC_1688 
+ TSMC_1689 TSMC_1690 TSMC_1691 TSMC_1692 TSMC_1693 TSMC_1694 
+ TSMC_1695 TSMC_1696 TSMC_1697 TSMC_1698 TSMC_1699 TSMC_1700 TSMC_1701 
+ TSMC_1702 TSMC_1703 TSMC_1704 TSMC_1705 TSMC_1706 TSMC_1707 
+ TSMC_1708 TSMC_1709 TSMC_1710 TSMC_1711 TSMC_1712 TSMC_1713 
+ TSMC_1714 TSMC_1715 TSMC_1716 TSMC_1717 TSMC_1718 TSMC_1719 
+ TSMC_1720 TSMC_1721 TSMC_1722 TSMC_1723 TSMC_1724 TSMC_1725 TSMC_1726 
+ TSMC_1727 TSMC_1728 TSMC_1729 TSMC_1730 TSMC_1731 TSMC_1732 
+ TSMC_1733 TSMC_1734 TSMC_1735 TSMC_1736 TSMC_1737 TSMC_1738 
+ TSMC_1739 TSMC_1740 TSMC_1741 TSMC_1742 TSMC_1743 TSMC_1744 TSMC_1745 
+ TSMC_1746 TSMC_1747 TSMC_1748 TSMC_1749 TSMC_1750 TSMC_1751 
+ TSMC_1752 TSMC_1753 TSMC_1754 TSMC_1755 TSMC_1756 TSMC_1757 
+ TSMC_1758 TSMC_1759 TSMC_1760 TSMC_1761 TSMC_1762 TSMC_1763 
+ S1ALLSVTSW2000X20_CELL_ARR_Y 
.ENDS

.SUBCKT S1ALLSVTSW2000X20_BOT_INOUT TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 
+ TSMC_7 TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 
+ TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 
+ TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 
+ TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 
+ TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 
+ TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 
+ TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 
+ TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 
+ TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 
+ TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 
+ TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 
+ TSMC_154 TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 
+ TSMC_162 TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 
+ TSMC_170 TSMC_171 TSMC_172 VDDHD VDDI TSMC_173 TSMC_174 VSSI TSMC_175 
+ TSMC_176 TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 
+ TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 
+ TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 
+ TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
XIO_L_0 TSMC_2 TSMC_34 TSMC_70 TSMC_103 TSMC_213 TSMC_135 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_1 TSMC_3 TSMC_35 TSMC_71 TSMC_104 TSMC_213 TSMC_136 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_2 TSMC_4 TSMC_36 TSMC_72 TSMC_105 TSMC_213 TSMC_137 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_3 TSMC_5 TSMC_37 TSMC_73 TSMC_106 TSMC_213 TSMC_138 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_4 TSMC_6 TSMC_38 TSMC_74 TSMC_107 TSMC_213 TSMC_139 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_5 TSMC_7 TSMC_39 TSMC_75 TSMC_108 TSMC_213 TSMC_140 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_6 TSMC_8 TSMC_40 TSMC_76 TSMC_109 TSMC_213 TSMC_141 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_7 TSMC_9 TSMC_41 TSMC_77 TSMC_110 TSMC_213 TSMC_142 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_8 TSMC_10 TSMC_42 TSMC_78 TSMC_111 TSMC_213 TSMC_143 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_9 TSMC_11 TSMC_43 TSMC_79 TSMC_112 TSMC_213 TSMC_144 VDDHD VDDI VSSI 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_10 TSMC_12 TSMC_44 TSMC_80 TSMC_113 TSMC_213 TSMC_145 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_11 TSMC_13 TSMC_45 TSMC_81 TSMC_114 TSMC_213 TSMC_146 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_12 TSMC_14 TSMC_46 TSMC_82 TSMC_115 TSMC_213 TSMC_147 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_L_13 TSMC_15 TSMC_47 TSMC_83 TSMC_116 TSMC_213 TSMC_148 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_18 TSMC_20 TSMC_52 TSMC_88 TSMC_121 TSMC_213 TSMC_153 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_19 TSMC_21 TSMC_53 TSMC_89 TSMC_122 TSMC_213 TSMC_154 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_20 TSMC_22 TSMC_54 TSMC_90 TSMC_123 TSMC_213 TSMC_155 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_21 TSMC_23 TSMC_55 TSMC_91 TSMC_124 TSMC_213 TSMC_156 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_22 TSMC_24 TSMC_56 TSMC_92 TSMC_125 TSMC_213 TSMC_157 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_23 TSMC_25 TSMC_57 TSMC_93 TSMC_126 TSMC_213 TSMC_158 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_24 TSMC_26 TSMC_58 TSMC_94 TSMC_127 TSMC_213 TSMC_159 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_25 TSMC_27 TSMC_59 TSMC_95 TSMC_128 TSMC_213 TSMC_160 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_26 TSMC_28 TSMC_60 TSMC_96 TSMC_129 TSMC_213 TSMC_161 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_27 TSMC_29 TSMC_61 TSMC_97 TSMC_130 TSMC_213 TSMC_162 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_28 TSMC_30 TSMC_62 TSMC_98 TSMC_131 TSMC_213 TSMC_163 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_29 TSMC_31 TSMC_63 TSMC_99 TSMC_132 TSMC_213 TSMC_164 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_30 TSMC_32 TSMC_64 TSMC_100 TSMC_133 TSMC_213 TSMC_165 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XIO_R_31 TSMC_33 TSMC_65 TSMC_101 TSMC_134 TSMC_213 TSMC_166 VDDHD VDDI 
+ VSSI S1ALLSVTSW2000X20_WOBIST_WOLS_IO_M8 
XCNTINOUT_M8 TSMC_1 TSMC_16 TSMC_19 TSMC_48 TSMC_51 TSMC_49 TSMC_50 
+ TSMC_17 TSMC_18 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_84 TSMC_87 TSMC_102 
+ TSMC_117 TSMC_120 TSMC_118 TSMC_119 TSMC_85 TSMC_86 TSMC_149 
+ TSMC_152 TSMC_150 TSMC_151 TSMC_167 TSMC_168 TSMC_174 TSMC_170 
+ TSMC_171 TSMC_172 VDDHD VDDI TSMC_173 TSMC_174 VSSI TSMC_175 TSMC_176 
+ TSMC_177 TSMC_178 TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 
+ TSMC_184 TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 
+ TSMC_191 TSMC_192 TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 
+ TSMC_199 TSMC_200 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ S1ALLSVTSW2000X20_WOBIST_WOLS_CNT_M8_IOX4 
.ENDS

.SUBCKT S1ALLSVTSW2000X20_BOT TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 
+ TSMC_8 TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_34 TSMC_35 
+ TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 
+ TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 
+ TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 
+ TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 
+ TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 
+ TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 
+ TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 
+ TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 
+ TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 TSMC_114 
+ TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 TSMC_122 
+ TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 
+ TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 
+ TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 
+ TSMC_147 TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 
+ TSMC_163 TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 
+ TSMC_171 TSMC_172 TSMC_173 TSMC_174 TSMC_175 TSMC_176 TSMC_177 TSMC_178 
+ TSMC_179 TSMC_180 TSMC_181 TSMC_182 TSMC_183 TSMC_184 TSMC_185 TSMC_186 
+ TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 TSMC_193 TSMC_194 
+ TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 TSMC_200 TSMC_201 TSMC_202 
+ TSMC_203 TSMC_204 TSMC_205 TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 
+ TSMC_211 TSMC_212 TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 
+ TSMC_219 TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 TSMC_234 
+ TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_239 TSMC_240 TSMC_241 TSMC_242 
+ TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_250 
+ TSMC_251 TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 
+ TSMC_259 TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 
+ TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_272 TSMC_273 TSMC_274 
+ TSMC_275 TSMC_276 TSMC_277 TSMC_278 TSMC_279 TSMC_280 TSMC_281 TSMC_282 
+ TSMC_283 TSMC_284 TSMC_285 TSMC_286 TSMC_287 TSMC_288 TSMC_289 TSMC_290 
+ TSMC_291 TSMC_292 TSMC_293 TSMC_294 TSMC_295 TSMC_296 TSMC_297 TSMC_298 
+ TSMC_299 TSMC_300 TSMC_301 VDDHD VDDI TSMC_302 TSMC_303 VSSI TSMC_304 
+ TSMC_305 TSMC_306 TSMC_307 TSMC_308 TSMC_309 TSMC_310 TSMC_311 TSMC_312 
+ TSMC_313 TSMC_314 TSMC_315 
XIO_L_0 TSMC_316 TSMC_18 TSMC_317 TSMC_95 TSMC_127 TSMC_159 TSMC_191 TSMC_223 
+ TSMC_318 TSMC_256 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_1 TSMC_316 TSMC_19 TSMC_317 TSMC_96 TSMC_128 TSMC_160 TSMC_192 TSMC_224 
+ TSMC_318 TSMC_257 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_2 TSMC_316 TSMC_20 TSMC_317 TSMC_97 TSMC_129 TSMC_161 TSMC_193 TSMC_225 
+ TSMC_318 TSMC_258 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_3 TSMC_316 TSMC_21 TSMC_317 TSMC_98 TSMC_130 TSMC_162 TSMC_194 TSMC_226 
+ TSMC_318 TSMC_259 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_4 TSMC_316 TSMC_22 TSMC_317 TSMC_99 TSMC_131 TSMC_163 TSMC_195 TSMC_227 
+ TSMC_318 TSMC_260 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_5 TSMC_316 TSMC_23 TSMC_317 TSMC_100 TSMC_132 TSMC_164 TSMC_196 TSMC_228 
+ TSMC_318 TSMC_261 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_6 TSMC_316 TSMC_24 TSMC_317 TSMC_101 TSMC_133 TSMC_165 TSMC_197 TSMC_229 
+ TSMC_318 TSMC_262 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_7 TSMC_316 TSMC_25 TSMC_317 TSMC_102 TSMC_134 TSMC_166 TSMC_198 TSMC_230 
+ TSMC_318 TSMC_263 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_8 TSMC_316 TSMC_26 TSMC_317 TSMC_103 TSMC_135 TSMC_167 TSMC_199 TSMC_231 
+ TSMC_318 TSMC_264 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_9 TSMC_316 TSMC_27 TSMC_317 TSMC_104 TSMC_136 TSMC_168 TSMC_200 TSMC_232 
+ TSMC_318 TSMC_265 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_10 TSMC_316 TSMC_28 TSMC_317 TSMC_105 TSMC_137 TSMC_169 TSMC_201 TSMC_233 
+ TSMC_318 TSMC_266 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_11 TSMC_316 TSMC_29 TSMC_317 TSMC_106 TSMC_138 TSMC_170 TSMC_202 TSMC_234 
+ TSMC_318 TSMC_267 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_12 TSMC_316 TSMC_30 TSMC_317 TSMC_107 TSMC_139 TSMC_171 TSMC_203 TSMC_235 
+ TSMC_318 TSMC_268 TSMC_319 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_L_13 TSMC_316 TSMC_31 TSMC_317 TSMC_108 TSMC_140 TSMC_172 TSMC_204 TSMC_236 
+ TSMC_322 TSMC_322 TSMC_318 TSMC_269 TSMC_296 TSMC_319 VDDHD VDDI 
+ VSSI TSMC_320 TSMC_321 S1ALLSVTSW2000X20_IO_M8 
XIO_R_18 TSMC_316 TSMC_36 TSMC_317 TSMC_113 TSMC_145 TSMC_177 TSMC_209 TSMC_241 
+ TSMC_322 TSMC_322 TSMC_323 TSMC_274 TSMC_296 TSMC_324 VDDHD VDDI 
+ VSSI TSMC_320 TSMC_321 S1ALLSVTSW2000X20_IO_M8 
XIO_R_19 TSMC_316 TSMC_37 TSMC_317 TSMC_114 TSMC_146 TSMC_178 TSMC_210 TSMC_242 
+ TSMC_323 TSMC_275 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_20 TSMC_316 TSMC_38 TSMC_317 TSMC_115 TSMC_147 TSMC_179 TSMC_211 TSMC_243 
+ TSMC_323 TSMC_276 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_21 TSMC_316 TSMC_39 TSMC_317 TSMC_116 TSMC_148 TSMC_180 TSMC_212 TSMC_244 
+ TSMC_323 TSMC_277 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_22 TSMC_316 TSMC_40 TSMC_317 TSMC_117 TSMC_149 TSMC_181 TSMC_213 TSMC_245 
+ TSMC_323 TSMC_278 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_23 TSMC_316 TSMC_41 TSMC_317 TSMC_118 TSMC_150 TSMC_182 TSMC_214 TSMC_246 
+ TSMC_323 TSMC_279 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_24 TSMC_316 TSMC_42 TSMC_317 TSMC_119 TSMC_151 TSMC_183 TSMC_215 TSMC_247 
+ TSMC_323 TSMC_280 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_25 TSMC_316 TSMC_43 TSMC_317 TSMC_120 TSMC_152 TSMC_184 TSMC_216 TSMC_248 
+ TSMC_323 TSMC_281 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_26 TSMC_316 TSMC_44 TSMC_317 TSMC_121 TSMC_153 TSMC_185 TSMC_217 TSMC_249 
+ TSMC_323 TSMC_282 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_27 TSMC_316 TSMC_45 TSMC_317 TSMC_122 TSMC_154 TSMC_186 TSMC_218 TSMC_250 
+ TSMC_323 TSMC_283 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_28 TSMC_316 TSMC_46 TSMC_317 TSMC_123 TSMC_155 TSMC_187 TSMC_219 TSMC_251 
+ TSMC_323 TSMC_284 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_29 TSMC_316 TSMC_47 TSMC_317 TSMC_124 TSMC_156 TSMC_188 TSMC_220 TSMC_252 
+ TSMC_323 TSMC_285 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_30 TSMC_316 TSMC_48 TSMC_317 TSMC_125 TSMC_157 TSMC_189 TSMC_221 TSMC_253 
+ TSMC_323 TSMC_286 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XIO_R_31 TSMC_316 TSMC_49 TSMC_317 TSMC_126 TSMC_158 TSMC_190 TSMC_222 TSMC_254 
+ TSMC_323 TSMC_287 TSMC_324 VDDHD VDDI VSSI TSMC_320 TSMC_321 
+ S1ALLSVTSW2000X20_IO_M8B 
XCNTIO_M8 TSMC_1 TSMC_316 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 
+ TSMC_9 TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 
+ TSMC_17 TSMC_32 TSMC_35 TSMC_33 TSMC_34 TSMC_50 TSMC_317 TSMC_51 
+ TSMC_51 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 TSMC_59 
+ TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 TSMC_67 
+ TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 TSMC_75 
+ TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 TSMC_83 
+ TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 TSMC_91 
+ TSMC_92 TSMC_93 TSMC_94 TSMC_109 TSMC_112 TSMC_110 TSMC_111 TSMC_141 
+ TSMC_144 TSMC_173 TSMC_176 TSMC_174 TSMC_175 TSMC_142 TSMC_143 
+ TSMC_205 TSMC_208 TSMC_237 TSMC_240 TSMC_238 TSMC_239 TSMC_206 TSMC_207 
+ TSMC_255 TSMC_325 TSMC_270 TSMC_273 TSMC_271 TSMC_272 TSMC_288 
+ TSMC_326 TSMC_327 TSMC_289 TSMC_290 TSMC_291 TSMC_292 TSMC_293 
+ TSMC_322 TSMC_322 TSMC_294 TSMC_296 TSMC_322 TSMC_295 TSMC_314 TSMC_315 
+ TSMC_328 TSMC_297 TSMC_298 TSMC_299 TSMC_300 TSMC_301 VDDHD VDDI 
+ TSMC_302 TSMC_303 VSSI TSMC_304 TSMC_305 TSMC_311 TSMC_306 TSMC_307 
+ TSMC_320 TSMC_308 TSMC_321 TSMC_309 TSMC_310 TSMC_312 TSMC_313 
+ S1ALLSVTSW2000X20_CNT_M8_IOX4 
.ENDS

.SUBCKT TS1N16FFCLLSVTA8192X32M8SW A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] A[8] 
+ A[9] A[10] A[11] A[12] BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] BWEB[5] 
+ BWEB[6] BWEB[7] BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12] BWEB[13] BWEB[14] 
+ BWEB[15] BWEB[16] BWEB[17] BWEB[18] BWEB[19] BWEB[20] BWEB[21] BWEB[22] 
+ BWEB[23] BWEB[24] BWEB[25] BWEB[26] BWEB[27] BWEB[28] BWEB[29] BWEB[30] 
+ BWEB[31] CEB CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] D[8] D[9] D[10] 
+ D[11] D[12] D[13] D[14] D[15] D[16] D[17] D[18] D[19] D[20] D[21] D[22] D[23] 
+ D[24] D[25] D[26] D[27] D[28] D[29] D[30] D[31] Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] 
+ Q[6] Q[7] Q[8] Q[9] Q[10] Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18] 
+ Q[19] Q[20] Q[21] Q[22] Q[23] Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] 
+ VDD VSS WEB WTSEL[0] WTSEL[1] RTSEL[0] RTSEL[1] 
XBANK0 TSMC_1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_24 TSMC_25 
+ TSMC_26 TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 
+ TSMC_34 TSMC_35 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 
+ TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 
+ TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 
+ TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 
+ TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 
+ TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 
+ TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 
+ TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 
+ TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 
+ TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 
+ TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 
+ TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 
+ TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 
+ TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 
+ TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 
+ TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 
+ TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 
+ TSMC_164 TSMC_165 TSMC_166 TSMC_167 TSMC_168 TSMC_169 TSMC_170 
+ TSMC_171 TSMC_172 VDD VDDHD VDD VSS TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ TSMC_177 TSMC_177 S1ALLSVTSW2000X20_BANK0_F 
XBANK1 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 TSMC_10 
+ TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 TSMC_18 
+ TSMC_19 TSMC_20 TSMC_21 TSMC_178 TSMC_179 TSMC_24 TSMC_25 TSMC_26 
+ TSMC_27 TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_32 TSMC_33 TSMC_35 
+ TSMC_180 TSMC_36 TSMC_37 TSMC_38 TSMC_39 TSMC_40 TSMC_41 TSMC_42 
+ TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 TSMC_48 TSMC_49 TSMC_50 
+ TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 TSMC_56 TSMC_57 TSMC_58 
+ TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 TSMC_64 TSMC_65 TSMC_66 
+ TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 TSMC_72 TSMC_73 TSMC_74 
+ TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 TSMC_80 TSMC_81 TSMC_82 
+ TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 TSMC_88 TSMC_89 TSMC_90 
+ TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 TSMC_96 TSMC_97 TSMC_98 TSMC_99 
+ TSMC_100 TSMC_101 TSMC_102 TSMC_103 TSMC_104 TSMC_105 TSMC_106 
+ TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 TSMC_112 TSMC_113 
+ TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 TSMC_119 TSMC_120 TSMC_121 
+ TSMC_122 TSMC_123 TSMC_124 TSMC_125 TSMC_126 TSMC_127 TSMC_128 
+ TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 TSMC_134 TSMC_135 
+ TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 TSMC_141 TSMC_142 TSMC_143 
+ TSMC_144 TSMC_145 TSMC_146 TSMC_147 TSMC_148 TSMC_149 TSMC_150 
+ TSMC_151 TSMC_152 TSMC_153 TSMC_154 TSMC_155 TSMC_156 TSMC_157 
+ TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 TSMC_163 TSMC_164 
+ TSMC_165 TSMC_167 TSMC_181 TSMC_182 TSMC_170 TSMC_183 TSMC_172 VDD 
+ VDDHD VDD VSS TSMC_173 TSMC_174 TSMC_175 TSMC_176 
+ S1ALLSVTSW2000X20_BANK_F 
XTOP_EDGE VDDHD VDD VSS TSMC_174 TSMC_184 S1ALLSVTSW2000X20_TOP_EDGE2 
XCNTIO TSMC_185 TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 TSMC_197 TSMC_198 TSMC_199 
+ TSMC_200 TSMC_1 TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 TSMC_233 CLK 
+ TSMC_234 TSMC_2 TSMC_3 TSMC_4 TSMC_5 TSMC_6 TSMC_7 TSMC_8 TSMC_9 
+ TSMC_10 TSMC_11 TSMC_12 TSMC_13 TSMC_14 TSMC_15 TSMC_16 TSMC_17 
+ TSMC_18 TSMC_19 TSMC_20 TSMC_21 TSMC_22 TSMC_23 TSMC_178 TSMC_179 
+ TSMC_235 TSMC_236 TSMC_237 TSMC_238 TSMC_24 TSMC_25 TSMC_26 TSMC_27 
+ TSMC_28 TSMC_29 TSMC_30 TSMC_31 TSMC_185 TSMC_32 TSMC_33 TSMC_239 
+ TSMC_239 TSMC_34 TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 
+ TSMC_245 TSMC_246 TSMC_247 TSMC_248 TSMC_249 TSMC_250 TSMC_251 
+ TSMC_252 TSMC_253 TSMC_254 TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 
+ TSMC_260 TSMC_261 TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 
+ TSMC_267 TSMC_268 TSMC_269 TSMC_270 TSMC_271 TSMC_36 TSMC_37 TSMC_38 
+ TSMC_39 TSMC_40 TSMC_41 TSMC_42 TSMC_43 TSMC_44 TSMC_45 TSMC_46 TSMC_47 
+ TSMC_48 TSMC_49 TSMC_50 TSMC_51 TSMC_52 TSMC_53 TSMC_54 TSMC_55 
+ TSMC_56 TSMC_57 TSMC_58 TSMC_59 TSMC_60 TSMC_61 TSMC_62 TSMC_63 
+ TSMC_64 TSMC_65 TSMC_66 TSMC_67 TSMC_68 TSMC_69 TSMC_70 TSMC_71 
+ TSMC_72 TSMC_73 TSMC_74 TSMC_75 TSMC_76 TSMC_77 TSMC_78 TSMC_79 
+ TSMC_80 TSMC_81 TSMC_82 TSMC_83 TSMC_84 TSMC_85 TSMC_86 TSMC_87 
+ TSMC_88 TSMC_89 TSMC_90 TSMC_91 TSMC_92 TSMC_93 TSMC_94 TSMC_95 
+ TSMC_96 TSMC_97 TSMC_98 TSMC_99 TSMC_100 TSMC_101 TSMC_102 TSMC_103 
+ TSMC_104 TSMC_105 TSMC_106 TSMC_107 TSMC_108 TSMC_109 TSMC_110 TSMC_111 
+ TSMC_112 TSMC_113 TSMC_114 TSMC_115 TSMC_116 TSMC_117 TSMC_118 
+ TSMC_119 TSMC_120 TSMC_121 TSMC_122 TSMC_123 TSMC_124 TSMC_125 
+ TSMC_126 TSMC_127 TSMC_128 TSMC_129 TSMC_130 TSMC_131 TSMC_132 TSMC_133 
+ TSMC_134 TSMC_135 TSMC_136 TSMC_137 TSMC_138 TSMC_139 TSMC_140 
+ TSMC_141 TSMC_142 TSMC_143 TSMC_144 TSMC_145 TSMC_146 TSMC_147 
+ TSMC_148 TSMC_149 TSMC_150 TSMC_151 TSMC_152 TSMC_153 TSMC_154 
+ TSMC_155 TSMC_156 TSMC_157 TSMC_158 TSMC_159 TSMC_160 TSMC_161 TSMC_162 
+ TSMC_163 TSMC_164 Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] 
+ Q[10] Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18] Q[19] Q[20] Q[21] 
+ Q[22] Q[23] Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] TSMC_165 
+ RTSEL[0] RTSEL[1] TSMC_185 TSMC_166 TSMC_182 TSMC_169 TSMC_185 
+ TSMC_272 TSMC_185 TSMC_185 TSMC_185 TSMC_172 TSMC_171 VDDHD VDD 
+ TSMC_239 TSMC_273 VSS TSMC_185 TSMC_185 TSMC_274 TSMC_174 TSMC_184 
+ WTSEL[0] WTSEL[1] TSMC_173 TSMC_175 TSMC_176 TSMC_177 TSMC_177 
+ S1ALLSVTSW2000X20_BOT 
XInput TSMC_185 BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] BWEB[5] BWEB[6] 
+ BWEB[7] BWEB[8] BWEB[9] BWEB[10] BWEB[11] BWEB[12] BWEB[13] BWEB[14] 
+ BWEB[15] BWEB[16] BWEB[17] BWEB[18] BWEB[19] BWEB[20] BWEB[21] BWEB[22] 
+ BWEB[23] BWEB[24] BWEB[25] BWEB[26] BWEB[27] BWEB[28] BWEB[29] 
+ BWEB[30] BWEB[31] TSMC_201 TSMC_202 TSMC_203 TSMC_204 TSMC_205 
+ TSMC_206 TSMC_207 TSMC_208 TSMC_209 TSMC_210 TSMC_211 TSMC_212 
+ TSMC_213 TSMC_214 TSMC_215 TSMC_216 TSMC_217 TSMC_218 TSMC_219 
+ TSMC_220 TSMC_221 TSMC_222 TSMC_223 TSMC_224 TSMC_225 TSMC_226 
+ TSMC_227 TSMC_228 TSMC_229 TSMC_230 TSMC_231 TSMC_232 CEB TSMC_233 
+ CLK TSMC_234 D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] D[8] D[9] D[10] 
+ D[11] D[12] D[13] D[14] D[15] D[16] D[17] D[18] D[19] D[20] D[21] D[22] 
+ D[23] D[24] D[25] D[26] D[27] D[28] D[29] D[30] D[31] TSMC_185 
+ TSMC_240 TSMC_241 TSMC_242 TSMC_243 TSMC_244 TSMC_245 TSMC_246 TSMC_247 
+ TSMC_248 TSMC_249 TSMC_250 TSMC_251 TSMC_252 TSMC_253 TSMC_254 
+ TSMC_255 TSMC_256 TSMC_257 TSMC_258 TSMC_259 TSMC_260 TSMC_261 
+ TSMC_262 TSMC_263 TSMC_264 TSMC_265 TSMC_266 TSMC_267 TSMC_268 TSMC_269 
+ TSMC_270 TSMC_271 Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] 
+ Q[10] Q[11] Q[12] Q[13] Q[14] Q[15] Q[16] Q[17] Q[18] Q[19] Q[20] Q[21] 
+ Q[22] Q[23] Q[24] Q[25] Q[26] Q[27] Q[28] Q[29] Q[30] Q[31] RTSEL[0] 
+ RTSEL[1] TSMC_185 TSMC_185 TSMC_185 TSMC_185 VDDHD VDD TSMC_275 
+ TSMC_185 VSS TSMC_185 TSMC_185 WEB TSMC_274 WTSEL[0] WTSEL[1] 
+ TSMC_186 TSMC_187 TSMC_188 TSMC_189 TSMC_190 TSMC_191 TSMC_192 
+ TSMC_193 TSMC_194 TSMC_195 TSMC_196 A[3] A[4] A[6] A[7] A[8] A[9] A[10] A[11] 
+ A[5] A[12] TSMC_185 TSMC_197 TSMC_198 TSMC_199 TSMC_200 A[0] A[1] A[2] 
+ TSMC_185 TSMC_177 TSMC_177 S1ALLSVTSW2000X20_BOT_INOUT 
XD_CEB CEB VSS S1ALLSVTSW2000X20_DIO 
XD_CLK CLK VSS S1ALLSVTSW2000X20_DIO 
XD_WEB WEB VSS S1ALLSVTSW2000X20_DIO 
XD_A0 A[0] VSS S1ALLSVTSW2000X20_DIO 
XD_A1 A[1] VSS S1ALLSVTSW2000X20_DIO 
XD_A2 A[2] VSS S1ALLSVTSW2000X20_DIO 
XD_A3 A[3] VSS S1ALLSVTSW2000X20_DIO 
XD_A4 A[4] VSS S1ALLSVTSW2000X20_DIO 
XD_A5 A[5] VSS S1ALLSVTSW2000X20_DIO 
XD_A6 A[6] VSS S1ALLSVTSW2000X20_DIO 
XD_A7 A[7] VSS S1ALLSVTSW2000X20_DIO 
XD_A8 A[8] VSS S1ALLSVTSW2000X20_DIO 
XD_A9 A[9] VSS S1ALLSVTSW2000X20_DIO 
XD_A10 A[10] VSS S1ALLSVTSW2000X20_DIO 
XD_A11 A[11] VSS S1ALLSVTSW2000X20_DIO 
XD_A12 A[12] VSS S1ALLSVTSW2000X20_DIO 
XD_D0 D[0] VSS S1ALLSVTSW2000X20_DIO 
XD_D1 D[1] VSS S1ALLSVTSW2000X20_DIO 
XD_D2 D[2] VSS S1ALLSVTSW2000X20_DIO 
XD_D3 D[3] VSS S1ALLSVTSW2000X20_DIO 
XD_D4 D[4] VSS S1ALLSVTSW2000X20_DIO 
XD_D5 D[5] VSS S1ALLSVTSW2000X20_DIO 
XD_D6 D[6] VSS S1ALLSVTSW2000X20_DIO 
XD_D7 D[7] VSS S1ALLSVTSW2000X20_DIO 
XD_D8 D[8] VSS S1ALLSVTSW2000X20_DIO 
XD_D9 D[9] VSS S1ALLSVTSW2000X20_DIO 
XD_D10 D[10] VSS S1ALLSVTSW2000X20_DIO 
XD_D11 D[11] VSS S1ALLSVTSW2000X20_DIO 
XD_D12 D[12] VSS S1ALLSVTSW2000X20_DIO 
XD_D13 D[13] VSS S1ALLSVTSW2000X20_DIO 
XD_D14 D[14] VSS S1ALLSVTSW2000X20_DIO 
XD_D15 D[15] VSS S1ALLSVTSW2000X20_DIO 
XD_D16 D[16] VSS S1ALLSVTSW2000X20_DIO 
XD_D17 D[17] VSS S1ALLSVTSW2000X20_DIO 
XD_D18 D[18] VSS S1ALLSVTSW2000X20_DIO 
XD_D19 D[19] VSS S1ALLSVTSW2000X20_DIO 
XD_D20 D[20] VSS S1ALLSVTSW2000X20_DIO 
XD_D21 D[21] VSS S1ALLSVTSW2000X20_DIO 
XD_D22 D[22] VSS S1ALLSVTSW2000X20_DIO 
XD_D23 D[23] VSS S1ALLSVTSW2000X20_DIO 
XD_D24 D[24] VSS S1ALLSVTSW2000X20_DIO 
XD_D25 D[25] VSS S1ALLSVTSW2000X20_DIO 
XD_D26 D[26] VSS S1ALLSVTSW2000X20_DIO 
XD_D27 D[27] VSS S1ALLSVTSW2000X20_DIO 
XD_D28 D[28] VSS S1ALLSVTSW2000X20_DIO 
XD_D29 D[29] VSS S1ALLSVTSW2000X20_DIO 
XD_D30 D[30] VSS S1ALLSVTSW2000X20_DIO 
XD_D31 D[31] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB0 BWEB[0] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB1 BWEB[1] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB2 BWEB[2] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB3 BWEB[3] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB4 BWEB[4] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB5 BWEB[5] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB6 BWEB[6] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB7 BWEB[7] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB8 BWEB[8] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB9 BWEB[9] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB10 BWEB[10] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB11 BWEB[11] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB12 BWEB[12] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB13 BWEB[13] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB14 BWEB[14] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB15 BWEB[15] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB16 BWEB[16] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB17 BWEB[17] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB18 BWEB[18] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB19 BWEB[19] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB20 BWEB[20] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB21 BWEB[21] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB22 BWEB[22] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB23 BWEB[23] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB24 BWEB[24] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB25 BWEB[25] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB26 BWEB[26] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB27 BWEB[27] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB28 BWEB[28] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB29 BWEB[29] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB30 BWEB[30] VSS S1ALLSVTSW2000X20_DIO 
XD_BWEB31 BWEB[31] VSS S1ALLSVTSW2000X20_DIO 
XD_WTSEL_1 WTSEL[1] VSS S1ALLSVTSW2000X20_DIO 
XD_WTSEL_0 WTSEL[0] VSS S1ALLSVTSW2000X20_DIO 
XD_RTSEL_1 RTSEL[1] VSS S1ALLSVTSW2000X20_DIO 
XD_RTSEL_0 RTSEL[0] VSS S1ALLSVTSW2000X20_DIO 
.ENDS


