# Created by MC2 : Version 2013.12.00.f on 2025/06/18, 13:11:27

 
###############################################################################
#                                                    
#        Technology     : TSMC 16nm CMOS Logic FinFet (FFC) HKMG
#        Memory Type    : TSMC 16nm FFC Two Port Register File with d130 bit cell
#        Library Name   : ts6n16ffcllsvta8x32m1fw (user specify : ts6n16ffcllsvta8x32m1fw)
#        Library Version: 170a
#        Generated Time : 2025/06/18, 13:10:29
###############################################################################
# STATEMENT OF USE                                                             
#                                                                              
#  This information contains confidential and proprietary information of TSMC. 
# No part of this information may be reproduced, transmitted, transcribed,     
# stored in a retrieval system, or translated into any human or computer       
# language, in any form or by any means, electronic, mechanical, magnetic,     
# optical, chemical, manual, or otherwise, without the prior written permission
# of TSMC. This information was prepared for informational purpose and is for  
# use by TSMC's customers only. TSMC reserves the right to make changes in the 
# inforrmation at any time and without notice.                                 
###############################################################################
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
#                                                                              

MACRO TS6N16FFCLLSVTA8X32M1FW
	CLASS BLOCK ;
	FOREIGN TS6N16FFCLLSVTA8X32M1FW 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 19.117 BY 43.680 ;
	SYMMETRY X Y ;
	PIN AA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 20.774 19.117 20.854 ;
			LAYER M2 ;
			RECT 18.869 20.774 19.117 20.854 ;
			LAYER M3 ;
			RECT 18.869 20.774 19.117 20.854 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[0]

	PIN AA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 19.178 19.117 19.258 ;
			LAYER M2 ;
			RECT 18.869 19.178 19.117 19.258 ;
			LAYER M3 ;
			RECT 18.869 19.178 19.117 19.258 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[1]

	PIN AA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 20.546 19.117 20.626 ;
			LAYER M2 ;
			RECT 18.869 20.546 19.117 20.626 ;
			LAYER M3 ;
			RECT 18.869 20.546 19.117 20.626 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0972 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2538 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AA[2]

	PIN AB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 22.826 19.117 22.906 ;
			LAYER M2 ;
			RECT 18.869 22.826 19.117 22.906 ;
			LAYER M3 ;
			RECT 18.869 22.826 19.117 22.906 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[0]

	PIN AB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 24.422 19.117 24.502 ;
			LAYER M2 ;
			RECT 18.869 24.422 19.117 24.502 ;
			LAYER M3 ;
			RECT 18.869 24.422 19.117 24.502 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[1]

	PIN AB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 23.054 19.117 23.134 ;
			LAYER M2 ;
			RECT 18.869 23.054 19.117 23.134 ;
			LAYER M3 ;
			RECT 18.869 23.054 19.117 23.134 ;
		END
		ANTENNAGATEAREA 0.0042 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0970 LAYER M1 ;
		ANTENNAMAXAREACAR 10.2024 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.2415 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0042 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1117 LAYER M2 ;
		ANTENNAMAXAREACAR 20.3208 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.4830 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0042 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5480 LAYER M3 ;
		ANTENNAMAXAREACAR 135.4520 LAYER M3 ;
	END AB[2]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 1.544 19.117 1.624 ;
			LAYER M2 ;
			RECT 18.869 1.544 19.117 1.624 ;
			LAYER M3 ;
			RECT 18.869 1.544 19.117 1.624 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 1.784 19.117 1.864 ;
			LAYER M2 ;
			RECT 18.869 1.784 19.117 1.864 ;
			LAYER M3 ;
			RECT 18.869 1.784 19.117 1.864 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 2.984 19.117 3.064 ;
			LAYER M2 ;
			RECT 18.869 2.984 19.117 3.064 ;
			LAYER M3 ;
			RECT 18.869 2.984 19.117 3.064 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 3.224 19.117 3.304 ;
			LAYER M2 ;
			RECT 18.869 3.224 19.117 3.304 ;
			LAYER M3 ;
			RECT 18.869 3.224 19.117 3.304 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 4.424 19.117 4.504 ;
			LAYER M2 ;
			RECT 18.869 4.424 19.117 4.504 ;
			LAYER M3 ;
			RECT 18.869 4.424 19.117 4.504 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 4.664 19.117 4.744 ;
			LAYER M2 ;
			RECT 18.869 4.664 19.117 4.744 ;
			LAYER M3 ;
			RECT 18.869 4.664 19.117 4.744 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 5.864 19.117 5.944 ;
			LAYER M2 ;
			RECT 18.869 5.864 19.117 5.944 ;
			LAYER M3 ;
			RECT 18.869 5.864 19.117 5.944 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 6.104 19.117 6.184 ;
			LAYER M2 ;
			RECT 18.869 6.104 19.117 6.184 ;
			LAYER M3 ;
			RECT 18.869 6.104 19.117 6.184 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 7.304 19.117 7.384 ;
			LAYER M2 ;
			RECT 18.869 7.304 19.117 7.384 ;
			LAYER M3 ;
			RECT 18.869 7.304 19.117 7.384 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 7.544 19.117 7.624 ;
			LAYER M2 ;
			RECT 18.869 7.544 19.117 7.624 ;
			LAYER M3 ;
			RECT 18.869 7.544 19.117 7.624 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[9]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 8.744 19.117 8.824 ;
			LAYER M2 ;
			RECT 18.869 8.744 19.117 8.824 ;
			LAYER M3 ;
			RECT 18.869 8.744 19.117 8.824 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 8.984 19.117 9.064 ;
			LAYER M2 ;
			RECT 18.869 8.984 19.117 9.064 ;
			LAYER M3 ;
			RECT 18.869 8.984 19.117 9.064 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 10.184 19.117 10.264 ;
			LAYER M2 ;
			RECT 18.869 10.184 19.117 10.264 ;
			LAYER M3 ;
			RECT 18.869 10.184 19.117 10.264 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 10.424 19.117 10.504 ;
			LAYER M2 ;
			RECT 18.869 10.424 19.117 10.504 ;
			LAYER M3 ;
			RECT 18.869 10.424 19.117 10.504 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 11.624 19.117 11.704 ;
			LAYER M2 ;
			RECT 18.869 11.624 19.117 11.704 ;
			LAYER M3 ;
			RECT 18.869 11.624 19.117 11.704 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 11.864 19.117 11.944 ;
			LAYER M2 ;
			RECT 18.869 11.864 19.117 11.944 ;
			LAYER M3 ;
			RECT 18.869 11.864 19.117 11.944 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 31.736 19.117 31.816 ;
			LAYER M2 ;
			RECT 18.869 31.736 19.117 31.816 ;
			LAYER M3 ;
			RECT 18.869 31.736 19.117 31.816 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 31.976 19.117 32.056 ;
			LAYER M2 ;
			RECT 18.869 31.976 19.117 32.056 ;
			LAYER M3 ;
			RECT 18.869 31.976 19.117 32.056 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 33.176 19.117 33.256 ;
			LAYER M2 ;
			RECT 18.869 33.176 19.117 33.256 ;
			LAYER M3 ;
			RECT 18.869 33.176 19.117 33.256 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 33.416 19.117 33.496 ;
			LAYER M2 ;
			RECT 18.869 33.416 19.117 33.496 ;
			LAYER M3 ;
			RECT 18.869 33.416 19.117 33.496 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 34.616 19.117 34.696 ;
			LAYER M2 ;
			RECT 18.869 34.616 19.117 34.696 ;
			LAYER M3 ;
			RECT 18.869 34.616 19.117 34.696 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 34.856 19.117 34.936 ;
			LAYER M2 ;
			RECT 18.869 34.856 19.117 34.936 ;
			LAYER M3 ;
			RECT 18.869 34.856 19.117 34.936 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 36.056 19.117 36.136 ;
			LAYER M2 ;
			RECT 18.869 36.056 19.117 36.136 ;
			LAYER M3 ;
			RECT 18.869 36.056 19.117 36.136 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 36.296 19.117 36.376 ;
			LAYER M2 ;
			RECT 18.869 36.296 19.117 36.376 ;
			LAYER M3 ;
			RECT 18.869 36.296 19.117 36.376 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 37.496 19.117 37.576 ;
			LAYER M2 ;
			RECT 18.869 37.496 19.117 37.576 ;
			LAYER M3 ;
			RECT 18.869 37.496 19.117 37.576 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 37.736 19.117 37.816 ;
			LAYER M2 ;
			RECT 18.869 37.736 19.117 37.816 ;
			LAYER M3 ;
			RECT 18.869 37.736 19.117 37.816 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 38.936 19.117 39.016 ;
			LAYER M2 ;
			RECT 18.869 38.936 19.117 39.016 ;
			LAYER M3 ;
			RECT 18.869 38.936 19.117 39.016 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 39.176 19.117 39.256 ;
			LAYER M2 ;
			RECT 18.869 39.176 19.117 39.256 ;
			LAYER M3 ;
			RECT 18.869 39.176 19.117 39.256 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 40.376 19.117 40.456 ;
			LAYER M2 ;
			RECT 18.869 40.376 19.117 40.456 ;
			LAYER M3 ;
			RECT 18.869 40.376 19.117 40.456 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 40.616 19.117 40.696 ;
			LAYER M2 ;
			RECT 18.869 40.616 19.117 40.696 ;
			LAYER M3 ;
			RECT 18.869 40.616 19.117 40.696 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 41.816 19.117 41.896 ;
			LAYER M2 ;
			RECT 18.869 41.816 19.117 41.896 ;
			LAYER M3 ;
			RECT 18.869 41.816 19.117 41.896 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 42.056 19.117 42.136 ;
			LAYER M2 ;
			RECT 18.869 42.056 19.117 42.136 ;
			LAYER M3 ;
			RECT 18.869 42.056 19.117 42.136 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2682 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3386 LAYER M3 ;
		ANTENNAMAXAREACAR 161.1170 LAYER M3 ;
	END BWEB[31]

	PIN CLKR
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 28.754 19.117 28.834 ;
			LAYER M2 ;
			RECT 18.869 28.754 19.117 28.834 ;
			LAYER M3 ;
			RECT 18.869 28.754 19.117 28.834 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2280 LAYER M2 ;
		ANTENNAMAXAREACAR 40.1766 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0128 LAYER M3 ;
		ANTENNAMAXAREACAR 179.9160 LAYER M3 ;
	END CLKR

	PIN CLKW
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 14.162 19.117 14.242 ;
			LAYER M2 ;
			RECT 18.869 14.162 19.117 14.242 ;
			LAYER M3 ;
			RECT 18.869 14.162 19.117 14.242 ;
		END
		ANTENNAGATEAREA 0.0060 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1144 LAYER M1 ;
		ANTENNAMAXAREACAR 11.0791 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0060 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.4639 LAYER M2 ;
		ANTENNAMAXAREACAR 44.8112 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0082 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0060 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 1.0159 LAYER M3 ;
		ANTENNAMAXAREACAR 150.9920 LAYER M3 ;
	END CLKW

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 1.064 19.117 1.144 ;
			LAYER M2 ;
			RECT 18.869 1.064 19.117 1.144 ;
			LAYER M3 ;
			RECT 18.869 1.064 19.117 1.144 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 2.264 19.117 2.344 ;
			LAYER M2 ;
			RECT 18.869 2.264 19.117 2.344 ;
			LAYER M3 ;
			RECT 18.869 2.264 19.117 2.344 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 2.504 19.117 2.584 ;
			LAYER M2 ;
			RECT 18.869 2.504 19.117 2.584 ;
			LAYER M3 ;
			RECT 18.869 2.504 19.117 2.584 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 3.704 19.117 3.784 ;
			LAYER M2 ;
			RECT 18.869 3.704 19.117 3.784 ;
			LAYER M3 ;
			RECT 18.869 3.704 19.117 3.784 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 3.944 19.117 4.024 ;
			LAYER M2 ;
			RECT 18.869 3.944 19.117 4.024 ;
			LAYER M3 ;
			RECT 18.869 3.944 19.117 4.024 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 5.144 19.117 5.224 ;
			LAYER M2 ;
			RECT 18.869 5.144 19.117 5.224 ;
			LAYER M3 ;
			RECT 18.869 5.144 19.117 5.224 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 5.384 19.117 5.464 ;
			LAYER M2 ;
			RECT 18.869 5.384 19.117 5.464 ;
			LAYER M3 ;
			RECT 18.869 5.384 19.117 5.464 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 6.584 19.117 6.664 ;
			LAYER M2 ;
			RECT 18.869 6.584 19.117 6.664 ;
			LAYER M3 ;
			RECT 18.869 6.584 19.117 6.664 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 6.824 19.117 6.904 ;
			LAYER M2 ;
			RECT 18.869 6.824 19.117 6.904 ;
			LAYER M3 ;
			RECT 18.869 6.824 19.117 6.904 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 8.024 19.117 8.104 ;
			LAYER M2 ;
			RECT 18.869 8.024 19.117 8.104 ;
			LAYER M3 ;
			RECT 18.869 8.024 19.117 8.104 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[9]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 8.264 19.117 8.344 ;
			LAYER M2 ;
			RECT 18.869 8.264 19.117 8.344 ;
			LAYER M3 ;
			RECT 18.869 8.264 19.117 8.344 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 9.464 19.117 9.544 ;
			LAYER M2 ;
			RECT 18.869 9.464 19.117 9.544 ;
			LAYER M3 ;
			RECT 18.869 9.464 19.117 9.544 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 9.704 19.117 9.784 ;
			LAYER M2 ;
			RECT 18.869 9.704 19.117 9.784 ;
			LAYER M3 ;
			RECT 18.869 9.704 19.117 9.784 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 10.904 19.117 10.984 ;
			LAYER M2 ;
			RECT 18.869 10.904 19.117 10.984 ;
			LAYER M3 ;
			RECT 18.869 10.904 19.117 10.984 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 11.144 19.117 11.224 ;
			LAYER M2 ;
			RECT 18.869 11.144 19.117 11.224 ;
			LAYER M3 ;
			RECT 18.869 11.144 19.117 11.224 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 12.344 19.117 12.424 ;
			LAYER M2 ;
			RECT 18.869 12.344 19.117 12.424 ;
			LAYER M3 ;
			RECT 18.869 12.344 19.117 12.424 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 31.256 19.117 31.336 ;
			LAYER M2 ;
			RECT 18.869 31.256 19.117 31.336 ;
			LAYER M3 ;
			RECT 18.869 31.256 19.117 31.336 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 32.456 19.117 32.536 ;
			LAYER M2 ;
			RECT 18.869 32.456 19.117 32.536 ;
			LAYER M3 ;
			RECT 18.869 32.456 19.117 32.536 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 32.696 19.117 32.776 ;
			LAYER M2 ;
			RECT 18.869 32.696 19.117 32.776 ;
			LAYER M3 ;
			RECT 18.869 32.696 19.117 32.776 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 33.896 19.117 33.976 ;
			LAYER M2 ;
			RECT 18.869 33.896 19.117 33.976 ;
			LAYER M3 ;
			RECT 18.869 33.896 19.117 33.976 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[19]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 34.136 19.117 34.216 ;
			LAYER M2 ;
			RECT 18.869 34.136 19.117 34.216 ;
			LAYER M3 ;
			RECT 18.869 34.136 19.117 34.216 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 35.336 19.117 35.416 ;
			LAYER M2 ;
			RECT 18.869 35.336 19.117 35.416 ;
			LAYER M3 ;
			RECT 18.869 35.336 19.117 35.416 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 35.576 19.117 35.656 ;
			LAYER M2 ;
			RECT 18.869 35.576 19.117 35.656 ;
			LAYER M3 ;
			RECT 18.869 35.576 19.117 35.656 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 36.776 19.117 36.856 ;
			LAYER M2 ;
			RECT 18.869 36.776 19.117 36.856 ;
			LAYER M3 ;
			RECT 18.869 36.776 19.117 36.856 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 37.016 19.117 37.096 ;
			LAYER M2 ;
			RECT 18.869 37.016 19.117 37.096 ;
			LAYER M3 ;
			RECT 18.869 37.016 19.117 37.096 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 38.216 19.117 38.296 ;
			LAYER M2 ;
			RECT 18.869 38.216 19.117 38.296 ;
			LAYER M3 ;
			RECT 18.869 38.216 19.117 38.296 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 38.456 19.117 38.536 ;
			LAYER M2 ;
			RECT 18.869 38.456 19.117 38.536 ;
			LAYER M3 ;
			RECT 18.869 38.456 19.117 38.536 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 39.656 19.117 39.736 ;
			LAYER M2 ;
			RECT 18.869 39.656 19.117 39.736 ;
			LAYER M3 ;
			RECT 18.869 39.656 19.117 39.736 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 39.896 19.117 39.976 ;
			LAYER M2 ;
			RECT 18.869 39.896 19.117 39.976 ;
			LAYER M3 ;
			RECT 18.869 39.896 19.117 39.976 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 41.096 19.117 41.176 ;
			LAYER M2 ;
			RECT 18.869 41.096 19.117 41.176 ;
			LAYER M3 ;
			RECT 18.869 41.096 19.117 41.176 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[29]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 41.336 19.117 41.416 ;
			LAYER M2 ;
			RECT 18.869 41.336 19.117 41.416 ;
			LAYER M3 ;
			RECT 18.869 41.336 19.117 41.416 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 42.536 19.117 42.616 ;
			LAYER M2 ;
			RECT 18.869 42.536 19.117 42.616 ;
			LAYER M3 ;
			RECT 18.869 42.536 19.117 42.616 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1465 LAYER M1 ;
		ANTENNAMAXAREACAR 7.6238 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2686 LAYER M2 ;
		ANTENNAMAXAREACAR 48.3629 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.2887 LAYER M3 ;
		ANTENNAMAXAREACAR 137.1780 LAYER M3 ;
	END D[31]

	PIN KP[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 15.530 19.117 15.610 ;
			LAYER M2 ;
			RECT 18.869 15.530 19.117 15.610 ;
			LAYER M3 ;
			RECT 18.869 15.530 19.117 15.610 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[0]

	PIN KP[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 15.758 19.117 15.838 ;
			LAYER M2 ;
			RECT 18.869 15.758 19.117 15.838 ;
			LAYER M3 ;
			RECT 18.869 15.758 19.117 15.838 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[1]

	PIN KP[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 15.986 19.117 16.066 ;
			LAYER M2 ;
			RECT 18.869 15.986 19.117 16.066 ;
			LAYER M3 ;
			RECT 18.869 15.986 19.117 16.066 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1415 LAYER M1 ;
		ANTENNAMAXAREACAR 16.7172 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.2401 LAYER M2 ;
		ANTENNAMAXAREACAR 29.3724 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0072 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.8346 LAYER M3 ;
		ANTENNAMAXAREACAR 329.2980 LAYER M3 ;
	END KP[2]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 1.304 19.117 1.384 ;
			LAYER M2 ;
			RECT 18.869 1.304 19.117 1.384 ;
			LAYER M3 ;
			RECT 18.869 1.304 19.117 1.384 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 2.024 19.117 2.104 ;
			LAYER M2 ;
			RECT 18.869 2.024 19.117 2.104 ;
			LAYER M3 ;
			RECT 18.869 2.024 19.117 2.104 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 2.744 19.117 2.824 ;
			LAYER M2 ;
			RECT 18.869 2.744 19.117 2.824 ;
			LAYER M3 ;
			RECT 18.869 2.744 19.117 2.824 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 3.464 19.117 3.544 ;
			LAYER M2 ;
			RECT 18.869 3.464 19.117 3.544 ;
			LAYER M3 ;
			RECT 18.869 3.464 19.117 3.544 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 4.184 19.117 4.264 ;
			LAYER M2 ;
			RECT 18.869 4.184 19.117 4.264 ;
			LAYER M3 ;
			RECT 18.869 4.184 19.117 4.264 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 4.904 19.117 4.984 ;
			LAYER M2 ;
			RECT 18.869 4.904 19.117 4.984 ;
			LAYER M3 ;
			RECT 18.869 4.904 19.117 4.984 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 5.624 19.117 5.704 ;
			LAYER M2 ;
			RECT 18.869 5.624 19.117 5.704 ;
			LAYER M3 ;
			RECT 18.869 5.624 19.117 5.704 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 6.344 19.117 6.424 ;
			LAYER M2 ;
			RECT 18.869 6.344 19.117 6.424 ;
			LAYER M3 ;
			RECT 18.869 6.344 19.117 6.424 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 7.064 19.117 7.144 ;
			LAYER M2 ;
			RECT 18.869 7.064 19.117 7.144 ;
			LAYER M3 ;
			RECT 18.869 7.064 19.117 7.144 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 7.784 19.117 7.864 ;
			LAYER M2 ;
			RECT 18.869 7.784 19.117 7.864 ;
			LAYER M3 ;
			RECT 18.869 7.784 19.117 7.864 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[9]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 8.504 19.117 8.584 ;
			LAYER M2 ;
			RECT 18.869 8.504 19.117 8.584 ;
			LAYER M3 ;
			RECT 18.869 8.504 19.117 8.584 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 9.224 19.117 9.304 ;
			LAYER M2 ;
			RECT 18.869 9.224 19.117 9.304 ;
			LAYER M3 ;
			RECT 18.869 9.224 19.117 9.304 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 9.944 19.117 10.024 ;
			LAYER M2 ;
			RECT 18.869 9.944 19.117 10.024 ;
			LAYER M3 ;
			RECT 18.869 9.944 19.117 10.024 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 10.664 19.117 10.744 ;
			LAYER M2 ;
			RECT 18.869 10.664 19.117 10.744 ;
			LAYER M3 ;
			RECT 18.869 10.664 19.117 10.744 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 11.384 19.117 11.464 ;
			LAYER M2 ;
			RECT 18.869 11.384 19.117 11.464 ;
			LAYER M3 ;
			RECT 18.869 11.384 19.117 11.464 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 12.104 19.117 12.184 ;
			LAYER M2 ;
			RECT 18.869 12.104 19.117 12.184 ;
			LAYER M3 ;
			RECT 18.869 12.104 19.117 12.184 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 31.496 19.117 31.576 ;
			LAYER M2 ;
			RECT 18.869 31.496 19.117 31.576 ;
			LAYER M3 ;
			RECT 18.869 31.496 19.117 31.576 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 32.216 19.117 32.296 ;
			LAYER M2 ;
			RECT 18.869 32.216 19.117 32.296 ;
			LAYER M3 ;
			RECT 18.869 32.216 19.117 32.296 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 32.936 19.117 33.016 ;
			LAYER M2 ;
			RECT 18.869 32.936 19.117 33.016 ;
			LAYER M3 ;
			RECT 18.869 32.936 19.117 33.016 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 33.656 19.117 33.736 ;
			LAYER M2 ;
			RECT 18.869 33.656 19.117 33.736 ;
			LAYER M3 ;
			RECT 18.869 33.656 19.117 33.736 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[19]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 34.376 19.117 34.456 ;
			LAYER M2 ;
			RECT 18.869 34.376 19.117 34.456 ;
			LAYER M3 ;
			RECT 18.869 34.376 19.117 34.456 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 35.096 19.117 35.176 ;
			LAYER M2 ;
			RECT 18.869 35.096 19.117 35.176 ;
			LAYER M3 ;
			RECT 18.869 35.096 19.117 35.176 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 35.816 19.117 35.896 ;
			LAYER M2 ;
			RECT 18.869 35.816 19.117 35.896 ;
			LAYER M3 ;
			RECT 18.869 35.816 19.117 35.896 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 36.536 19.117 36.616 ;
			LAYER M2 ;
			RECT 18.869 36.536 19.117 36.616 ;
			LAYER M3 ;
			RECT 18.869 36.536 19.117 36.616 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 37.256 19.117 37.336 ;
			LAYER M2 ;
			RECT 18.869 37.256 19.117 37.336 ;
			LAYER M3 ;
			RECT 18.869 37.256 19.117 37.336 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 37.976 19.117 38.056 ;
			LAYER M2 ;
			RECT 18.869 37.976 19.117 38.056 ;
			LAYER M3 ;
			RECT 18.869 37.976 19.117 38.056 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 38.696 19.117 38.776 ;
			LAYER M2 ;
			RECT 18.869 38.696 19.117 38.776 ;
			LAYER M3 ;
			RECT 18.869 38.696 19.117 38.776 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 39.416 19.117 39.496 ;
			LAYER M2 ;
			RECT 18.869 39.416 19.117 39.496 ;
			LAYER M3 ;
			RECT 18.869 39.416 19.117 39.496 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 40.136 19.117 40.216 ;
			LAYER M2 ;
			RECT 18.869 40.136 19.117 40.216 ;
			LAYER M3 ;
			RECT 18.869 40.136 19.117 40.216 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 40.856 19.117 40.936 ;
			LAYER M2 ;
			RECT 18.869 40.856 19.117 40.936 ;
			LAYER M3 ;
			RECT 18.869 40.856 19.117 40.936 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[29]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 41.576 19.117 41.656 ;
			LAYER M2 ;
			RECT 18.869 41.576 19.117 41.656 ;
			LAYER M3 ;
			RECT 18.869 41.576 19.117 41.656 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 42.296 19.117 42.376 ;
			LAYER M2 ;
			RECT 18.869 42.296 19.117 42.376 ;
			LAYER M3 ;
			RECT 18.869 42.296 19.117 42.376 ;
		END
		ANTENNADIFFAREA 0.0566 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1328 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNADIFFAREA 0.0566 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1391 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNADIFFAREA 0.0566 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.3720 LAYER M3 ;
	END Q[31]

	PIN RCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 30.578 19.117 30.658 ;
			LAYER M2 ;
			RECT 18.869 30.578 19.117 30.658 ;
			LAYER M3 ;
			RECT 18.869 30.578 19.117 30.658 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[0]

	PIN RCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 30.350 19.117 30.430 ;
			LAYER M2 ;
			RECT 18.869 30.350 19.117 30.430 ;
			LAYER M3 ;
			RECT 18.869 30.350 19.117 30.430 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1188 LAYER M1 ;
		ANTENNAMAXAREACAR 17.6586 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1107 LAYER M2 ;
		ANTENNAMAXAREACAR 39.0207 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5592 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8850 LAYER M3 ;
	END RCT[1]

	PIN REB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 26.930 19.117 27.010 ;
			LAYER M2 ;
			RECT 18.869 26.930 19.117 27.010 ;
			LAYER M3 ;
			RECT 18.869 26.930 19.117 27.010 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0860 LAYER M1 ;
		ANTENNAMAXAREACAR 12.8828 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0840 LAYER M2 ;
		ANTENNAMAXAREACAR 20.5069 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4602 LAYER M3 ;
		ANTENNAMAXAREACAR 218.8550 LAYER M3 ;
	END REB

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.120 1.624 18.997 1.784 ;
			LAYER M4 ;
			RECT 0.120 3.064 18.997 3.224 ;
			LAYER M4 ;
			RECT 0.120 4.504 18.997 4.664 ;
			LAYER M4 ;
			RECT 0.120 5.944 18.997 6.104 ;
			LAYER M4 ;
			RECT 0.120 7.384 18.997 7.544 ;
			LAYER M4 ;
			RECT 0.120 8.824 18.997 8.984 ;
			LAYER M4 ;
			RECT 0.120 10.264 18.997 10.424 ;
			LAYER M4 ;
			RECT 0.120 11.704 18.997 11.864 ;
			LAYER M4 ;
			RECT 0.120 13.124 18.997 13.324 ;
			LAYER M4 ;
			RECT 0.120 14.060 18.997 14.260 ;
			LAYER M4 ;
			RECT 0.120 15.596 18.997 15.796 ;
			LAYER M4 ;
			RECT 0.120 17.132 18.997 17.332 ;
			LAYER M4 ;
			RECT 0.120 18.668 18.997 18.868 ;
			LAYER M4 ;
			RECT 0.120 20.204 18.997 20.404 ;
			LAYER M4 ;
			RECT 0.120 21.740 18.997 21.940 ;
			LAYER M4 ;
			RECT 0.120 23.276 18.997 23.476 ;
			LAYER M4 ;
			RECT 0.120 24.812 18.997 25.012 ;
			LAYER M4 ;
			RECT 0.120 26.348 18.997 26.548 ;
			LAYER M4 ;
			RECT 0.120 27.884 18.997 28.084 ;
			LAYER M4 ;
			RECT 0.120 29.420 18.997 29.620 ;
			LAYER M4 ;
			RECT 0.120 30.356 18.997 30.556 ;
			LAYER M4 ;
			RECT 0.120 31.816 18.997 31.976 ;
			LAYER M4 ;
			RECT 0.120 33.256 18.997 33.416 ;
			LAYER M4 ;
			RECT 0.120 34.696 18.997 34.856 ;
			LAYER M4 ;
			RECT 0.120 36.136 18.997 36.296 ;
			LAYER M4 ;
			RECT 0.120 37.576 18.997 37.736 ;
			LAYER M4 ;
			RECT 0.120 39.016 18.997 39.176 ;
			LAYER M4 ;
			RECT 0.120 40.456 18.997 40.616 ;
			LAYER M4 ;
			RECT 0.120 41.896 18.997 42.056 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.120 0.884 18.997 1.084 ;
			LAYER M4 ;
			RECT 0.120 2.324 18.997 2.524 ;
			LAYER M4 ;
			RECT 0.120 3.764 18.997 3.964 ;
			LAYER M4 ;
			RECT 0.120 5.204 18.997 5.404 ;
			LAYER M4 ;
			RECT 0.120 6.644 18.997 6.844 ;
			LAYER M4 ;
			RECT 0.120 8.084 18.997 8.284 ;
			LAYER M4 ;
			RECT 0.120 9.524 18.997 9.724 ;
			LAYER M4 ;
			RECT 0.120 10.964 18.997 11.164 ;
			LAYER M4 ;
			RECT 0.120 12.404 18.997 12.604 ;
			LAYER M4 ;
			RECT 0.120 14.828 18.997 15.028 ;
			LAYER M4 ;
			RECT 0.120 16.364 18.997 16.564 ;
			LAYER M4 ;
			RECT 0.120 17.900 18.997 18.100 ;
			LAYER M4 ;
			RECT 0.120 19.436 18.997 19.636 ;
			LAYER M4 ;
			RECT 0.120 20.972 18.997 21.172 ;
			LAYER M4 ;
			RECT 0.120 22.508 18.997 22.708 ;
			LAYER M4 ;
			RECT 0.120 24.044 18.997 24.244 ;
			LAYER M4 ;
			RECT 0.120 25.580 18.997 25.780 ;
			LAYER M4 ;
			RECT 0.120 27.116 18.997 27.316 ;
			LAYER M4 ;
			RECT 0.120 28.652 18.997 28.852 ;
			LAYER M4 ;
			RECT 0.120 31.076 18.997 31.276 ;
			LAYER M4 ;
			RECT 0.120 32.516 18.997 32.716 ;
			LAYER M4 ;
			RECT 0.120 33.956 18.997 34.156 ;
			LAYER M4 ;
			RECT 0.120 35.396 18.997 35.596 ;
			LAYER M4 ;
			RECT 0.120 36.836 18.997 37.036 ;
			LAYER M4 ;
			RECT 0.120 38.276 18.997 38.476 ;
			LAYER M4 ;
			RECT 0.120 39.716 18.997 39.916 ;
			LAYER M4 ;
			RECT 0.120 41.156 18.997 41.356 ;
			LAYER M4 ;
			RECT 0.120 42.596 18.997 42.796 ;
		END
	END VSS

	PIN WCT[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 13.478 19.117 13.558 ;
			LAYER M2 ;
			RECT 18.869 13.478 19.117 13.558 ;
			LAYER M3 ;
			RECT 18.869 13.478 19.117 13.558 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[0]

	PIN WCT[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 13.250 19.117 13.330 ;
			LAYER M2 ;
			RECT 18.869 13.250 19.117 13.330 ;
			LAYER M3 ;
			RECT 18.869 13.250 19.117 13.330 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.1482 LAYER M1 ;
		ANTENNAMAXAREACAR 16.9345 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.1043 LAYER M2 ;
		ANTENNAMAXAREACAR 44.5966 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0051 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.5855 LAYER M3 ;
		ANTENNAMAXAREACAR 105.8140 LAYER M3 ;
	END WCT[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.869 16.670 19.117 16.750 ;
			LAYER M2 ;
			RECT 18.869 16.670 19.117 16.750 ;
			LAYER M3 ;
			RECT 18.869 16.670 19.117 16.750 ;
		END
		ANTENNAGATEAREA 0.0023 LAYER M1 ;
		ANTENNADIFFAREA 0.0081 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.0886 LAYER M1 ;
		ANTENNAMAXAREACAR 9.6368 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.4414 LAYER VIA1 ;
		ANTENNAGATEAREA 0.0023 LAYER M2 ;
		ANTENNADIFFAREA 0.0081 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.0833 LAYER M2 ;
		ANTENNAMAXAREACAR 13.2425 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.0041 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.8828 LAYER VIA2 ;
		ANTENNAGATEAREA 0.0023 LAYER M3 ;
		ANTENNADIFFAREA 0.0081 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.4593 LAYER M3 ;
		ANTENNAMAXAREACAR 211.0720 LAYER M3 ;
	END WEB

	OBS
		LAYER M1 ;
		RECT 0.000 0.000 19.117 43.680 ;
		LAYER M2 ;
		RECT 0.000 0.000 19.117 43.680 ;
		LAYER M3 ;
		RECT 0.000 0.000 19.117 43.680 ;
		LAYER M4 ;
		RECT 0.227 0.524 18.567 0.724 ;
		LAYER M4 ;
		RECT 0.227 1.358 18.137 1.518 ;
		LAYER M4 ;
		RECT 0.227 1.890 18.137 2.050 ;
		LAYER M4 ;
		RECT 0.227 2.798 18.137 2.958 ;
		LAYER M4 ;
		RECT 0.227 3.330 18.137 3.490 ;
		LAYER M4 ;
		RECT 0.227 4.238 18.137 4.398 ;
		LAYER M4 ;
		RECT 0.227 4.770 18.137 4.930 ;
		LAYER M4 ;
		RECT 0.227 5.678 18.137 5.838 ;
		LAYER M4 ;
		RECT 0.227 6.210 18.137 6.370 ;
		LAYER M4 ;
		RECT 0.227 7.118 18.137 7.278 ;
		LAYER M4 ;
		RECT 0.227 7.650 18.137 7.810 ;
		LAYER M4 ;
		RECT 0.227 8.558 18.137 8.718 ;
		LAYER M4 ;
		RECT 0.227 9.090 18.137 9.250 ;
		LAYER M4 ;
		RECT 0.227 9.998 18.137 10.158 ;
		LAYER M4 ;
		RECT 0.227 10.530 18.137 10.690 ;
		LAYER M4 ;
		RECT 0.227 11.438 18.137 11.598 ;
		LAYER M4 ;
		RECT 0.227 11.970 18.137 12.130 ;
		LAYER M4 ;
		RECT 0.227 12.764 18.137 12.964 ;
		LAYER M4 ;
		RECT 0.227 13.676 18.137 13.876 ;
		LAYER M4 ;
		RECT 0.227 14.444 18.137 14.644 ;
		LAYER M4 ;
		RECT 0.227 15.212 18.137 15.412 ;
		LAYER M4 ;
		RECT 0.227 15.980 18.137 16.180 ;
		LAYER M4 ;
		RECT 0.227 16.748 18.137 16.948 ;
		LAYER M4 ;
		RECT 0.227 17.516 18.137 17.716 ;
		LAYER M4 ;
		RECT 0.227 18.284 18.137 18.484 ;
		LAYER M4 ;
		RECT 0.227 19.052 18.137 19.252 ;
		LAYER M4 ;
		RECT 0.227 19.820 18.137 20.020 ;
		LAYER M4 ;
		RECT 0.227 20.588 18.137 20.788 ;
		LAYER M4 ;
		RECT 0.227 21.356 18.137 21.556 ;
		LAYER M4 ;
		RECT 0.227 22.124 18.137 22.324 ;
		LAYER M4 ;
		RECT 0.227 22.892 18.137 23.092 ;
		LAYER M4 ;
		RECT 0.227 23.660 18.137 23.860 ;
		LAYER M4 ;
		RECT 0.227 24.428 18.137 24.628 ;
		LAYER M4 ;
		RECT 0.227 25.196 18.137 25.396 ;
		LAYER M4 ;
		RECT 0.227 25.964 18.137 26.164 ;
		LAYER M4 ;
		RECT 0.227 26.732 18.137 26.932 ;
		LAYER M4 ;
		RECT 0.227 27.500 18.137 27.700 ;
		LAYER M4 ;
		RECT 0.227 28.268 18.137 28.468 ;
		LAYER M4 ;
		RECT 0.227 29.036 18.137 29.236 ;
		LAYER M4 ;
		RECT 0.227 29.804 18.137 30.004 ;
		LAYER M4 ;
		RECT 0.227 30.716 18.137 30.916 ;
		LAYER M4 ;
		RECT 0.227 31.550 18.137 31.710 ;
		LAYER M4 ;
		RECT 0.227 32.082 18.137 32.242 ;
		LAYER M4 ;
		RECT 0.227 32.990 18.137 33.150 ;
		LAYER M4 ;
		RECT 0.227 33.522 18.137 33.682 ;
		LAYER M4 ;
		RECT 0.227 34.430 18.137 34.590 ;
		LAYER M4 ;
		RECT 0.227 34.962 18.137 35.122 ;
		LAYER M4 ;
		RECT 0.227 35.870 18.137 36.030 ;
		LAYER M4 ;
		RECT 0.227 36.402 18.137 36.562 ;
		LAYER M4 ;
		RECT 0.227 37.310 18.137 37.470 ;
		LAYER M4 ;
		RECT 0.227 37.842 18.137 38.002 ;
		LAYER M4 ;
		RECT 0.227 38.750 18.137 38.910 ;
		LAYER M4 ;
		RECT 0.227 39.282 18.137 39.442 ;
		LAYER M4 ;
		RECT 0.227 40.190 18.137 40.350 ;
		LAYER M4 ;
		RECT 0.227 40.722 18.137 40.882 ;
		LAYER M4 ;
		RECT 0.227 41.630 18.137 41.790 ;
		LAYER M4 ;
		RECT 0.227 42.162 18.137 42.322 ;
		LAYER M4 ;
		RECT 0.227 42.956 18.567 43.156 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 19.117 43.680 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 19.117 43.680 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 19.117 43.680 ;
	END
END TS6N16FFCLLSVTA8X32M1FW

END LIBRARY
